/*
date:2018/5/8
���ںţ�С��FPGA
���ں��ϡ���2Ƶ��FFTʵ��-verilogƪ2�������̽���
*/

module fw_sram_1 #(
  parameter WIDTH_A = 12
)
(
   input [WIDTH_A-1:0] addr,
   
   output[119:0]  coef

);

       

wire [119:0] Coef [0:1273];
assign Coef[0] = 'hFF5B6BD14C3E55E340906C1DEB5F67;
assign Coef[1] = 'hD1EB735A4DE679C30B95BF2DC09E77;
assign Coef[2] = 'hF76248CADE083F81C1B6E9AF925C61;
assign Coef[3] = 'hF5C05B4A6C802D6261B0D8FE9B17E9;
assign Coef[4] = 'h457656484E20AD63F7B4BAD7951DD1;
assign Coef[5] = 'h5F5BCAC846863D6346D27C3FDA19E7;
assign Coef[6] = 'hAE17F949C722B523775950BF97B26B;
assign Coef[7] = 'h486BEED134254E76F7E8626BF52FBC;
assign Coef[8] = 'h96DD59BA21C7BCCDF5B3668E543292;
assign Coef[9] = 'h2620F89A3775BB55705A76ED04EA35;
assign Coef[10] = 'hAE21AA01524FA47D7746DE9AA0E0BC;
assign Coef[11] = 'hB8357B92104F3ACB3402070C085D02;
assign Coef[12] = 'hA9EB18DA63F269617098B406B57990;
assign Coef[13] = 'hB72151C06CEC752B05EA33AF72D564;
assign Coef[14] = 'h2D7F42F35D1C38EB451C697B85C66D;
assign Coef[15] = 'h29700DC269349B82A3B2081B439045;
assign Coef[16] = 'hEA5C5008492067E342BEE474E89A6C;
assign Coef[17] = 'h1F4A9CF85CACE34277EE898AF71200;
assign Coef[18] = 'hBB8A7243AE94216A7061E20B7284C1;
assign Coef[19] = 'h802FEA4344BD66D362FDD6CA9E2295;
assign Coef[20] = 'h936D39A90337E64962F2F2F8EAF121;
assign Coef[21] = 'h525D7F91305FD2D5777A76ECA2F138;
assign Coef[22] = 'h2258FCB1B117405E97FAC47883F102;
assign Coef[23] = 'h8A8DE3A9224FFEFF6DC77A68047B12;
assign Coef[24] = 'h06097FB0225BFE7766DF64CC917310;
assign Coef[25] = 'h0ADD78B9318FE2B7F5CE4069637A0A;
assign Coef[26] = 'hDD1A77F35C1CF7476099BCD8F18EED;
assign Coef[27] = 'hC5FB6848CE2C15C6B182F809AB9DF9;
assign Coef[28] = 'hE1E24B635CAC3560F18BFD8FB60CE9;
assign Coef[29] = 'hDD7AD1504C8021A3B79402BB7391E9;
assign Coef[30] = 'hD575424A9BA089E3C3A6FAEE2C05F9;
assign Coef[31] = 'hD7D253417FAC22E35383945E7199DC;
assign Coef[32] = 'hCFE15A9A25C28DC557F4209E553F12;
assign Coef[33] = 'h893B48987787F143C3D7585B05BF83;
assign Coef[34] = 'h3651FDB82167B3D767657C4143F83A;
assign Coef[35] = 'hAC1554B8E15DE0D5E61E541D41F736;
assign Coef[36] = 'h0858C3B333DFEDD7F050D4D984EB36;
assign Coef[37] = 'h1EBA7FB9605E3156039262E171FAE7;
assign Coef[38] = 'h7695C1194C12B04022C3B21239716B;
assign Coef[39] = 'hA3B3534366C4AB619175662F5ECDE4;
assign Coef[40] = 'hFF36D8F08C94726345F2923D54956D;
assign Coef[41] = 'h625A43DB7DA075662064F67E0352ED;
assign Coef[42] = 'h63BB6173CDE02467DC1EEF0E33814A;
assign Coef[43] = 'h7DCB5F6BA20C6D41EC2F3749948EED;
assign Coef[44] = 'hE5DC69CB7C443749653F60989383D7;
assign Coef[45] = 'hF239F4FA66D566A792B6D220E7B6B2;
assign Coef[46] = 'hE2CECCAB12DEBF65F1EB9009BDBAE9;
assign Coef[47] = 'h9071E320E35D6486236F742DA5F15A;
assign Coef[48] = 'h1AD97EBA7277E075573C52ADA5EB36;
assign Coef[49] = 'h88C9F631237D93F7075904F823EA8C;
assign Coef[50] = 'h08E9A03030FFE2D6F74166E02F6218;
assign Coef[51] = 'h1A5D77B1A37FAAC7D7504648B5FF8C;
assign Coef[52] = 'h81CB27715C7EB605610329EDE72F32;
assign Coef[53] = 'hD1FA51531D0871A171932DEC799AD9;
assign Coef[54] = 'hF5CAD34ADEE87DC2B0AFF5CC738E75;
assign Coef[55] = 'hD77341D34A445F41F09ADEAF56DE73;
assign Coef[56] = 'hF6D20D43A896B0C79196F04F788CEA;
assign Coef[57] = 'h7127D47327A4094155E2E8DBC4B5AE;
assign Coef[58] = 'h4F6F7FF837AD222BF7B758CB02A4BC;
assign Coef[59] = 'h589DE59230EFBB6AC6587A3345FA82;
assign Coef[60] = 'h08FD469233D7B78457E96E8935F49E;
assign Coef[61] = 'h48F86DB1B3D7A9B5F7406641456FBF;
assign Coef[62] = 'h2A1F4D3BB1F779DF41D8140B25F8C6;
assign Coef[63] = 'h267C5539664FF22143C77E2C6C983C;
assign Coef[64] = 'h0E77560040B6340304D8B81BC1BD0F;
assign Coef[65] = 'h3BE95D52039447F003F44A3F2E55FC;
assign Coef[66] = 'hE4755E4BFD302C45104BE4CE44941F;
assign Coef[67] = 'h65FFD9CACE966F61300C0ECF57C737;
assign Coef[68] = 'hB6E312280C9CA5A2809B6E4EDD8B69;
assign Coef[69] = 'hEB66D06B8F9C7FC5E4A0B96BC383F2;
assign Coef[70] = 'hCF4B566B480743806DBA6B9BB28EE1;
assign Coef[71] = 'h030AD6421696CE412029507F17CD54;
assign Coef[72] = 'h36024029F7632BC0266DF56810D8A9;
assign Coef[73] = 'hAE2DF520B95F52E5D5627E7FE7E133;
assign Coef[74] = 'h6E89E5A020D5B7F735452BAE64F0BC;
assign Coef[75] = 'h5C49742163DFE89367DD34ECE2EFAC;
assign Coef[76] = 'hDA0964B1B2FFEE75136F40C8E9E08C;
assign Coef[77] = 'h2899072973D7E7A6F7E26219A1FB1A;
assign Coef[78] = 'hA74A57792EC67061A39A3E5F21CFDD;
assign Coef[79] = 'h33520A6ACC0431C1F08F3E8BD095C9;
assign Coef[80] = 'hC56348FA4EA87BE8D982BD8FC4066D;
assign Coef[81] = 'h7477187A4700166C2181EE9F77C77A;
assign Coef[82] = 'hC07E00D86C0025C5E13F48DCD00C19;
assign Coef[83] = 'h7A230C0BD50138E1F7380A56559CC2;
assign Coef[84] = 'h4815088825816A629513228C17FE96;
assign Coef[85] = 'h14705F9A11EFE557E5DB6889E62F84;
assign Coef[86] = 'h2AD4089333C3F875C65048C138FAB6;
assign Coef[87] = 'h52501EACB177DA3507641E5D6075F7;
assign Coef[88] = 'h0829C0B922FFB2CD31D368717FE514;
assign Coef[89] = 'hBAB8DDB923FD7E8110F31C3B26F226;
assign Coef[90] = 'h75E406D3778EE8C7016A6EFA9E9B73;
assign Coef[91] = 'h642200C207B7EA0D8392F07E3E96A1;
assign Coef[92] = 'hDFE754F975243D0B15FE3EADD3037D;
assign Coef[93] = 'h7D1246714C0229A156AC3DCFD253E4;
assign Coef[94] = 'h2DB550484C6075C722A75CAF8BC76D;
assign Coef[95] = 'h77BC52437E9F119246A7792EF78763;
assign Coef[96] = 'hB3134A424EF5F857B74152D6DF9684;
assign Coef[97] = 'h325B490AEA15BE53161E6288EAD8C7;
assign Coef[98] = 'h18095C40E1679B47A7DD56152BB05C;
assign Coef[99] = 'h10894CB02366ECC793E6286826327C;
assign Coef[100] = 'h62C98CA12117AE6012E128E914EB2A;
assign Coef[101] = 'h5ADD4AA8326FF864E6F860682DFA1B;
assign Coef[102] = 'h2695D6A1227F6370E3C646C800F90A;
assign Coef[103] = 'h4C8D9EA0A3FF6587156D24E8F7A9BE;
assign Coef[104] = 'hD1050E702C56CD85F19FADDFA28468;
assign Coef[105] = 'h612B507ECF741B03E896ACCBD69571;
assign Coef[106] = 'hA572C0FACF9829E0B88DBEFF5256E4;
assign Coef[107] = 'h737142EBD54448C3E719B89F72557D;
assign Coef[108] = 'h837442C954068CA2A0B168FF741667;
assign Coef[109] = 'h4C771202412042D129AC3C9F7284F2;
assign Coef[110] = 'h0E648791716ED4674F3F3E6A157C0B;
assign Coef[111] = 'hDA799F96A1C7DFF135160A7C612E1F;
assign Coef[112] = 'h4E78379E31D3BC7C23F31E11C5EA8E;
assign Coef[113] = 'h187CCBB1A1DFEC9637F02ED880EA13;
assign Coef[114] = 'h582CD13F31DFBA7D134E6E0B5CFB37;
assign Coef[115] = 'h3E24D03753CABD23017F7C7CD08B02;
assign Coef[116] = 'h64740A08A5240D05EA713CB821F4E1;
assign Coef[117] = 'h6762124141048F2B91A5721DFC94D0;
assign Coef[118] = 'h4F3846525E1038A0022EFA0E3606CE;
assign Coef[119] = 'h633ECE386F94288190A7050E1602ED;
assign Coef[120] = 'h1F880EB0ECA466C10C133D0F120775;
assign Coef[121] = 'hCDE248A91F840D42B21649AE9E8DC9;
assign Coef[122] = 'hC31E456C059C294777A26A2E210508;
assign Coef[123] = 'h8F0F938E96457DF1A62E2CAC013F32;
assign Coef[124] = 'h7219C4A11755E84595A918040222F7;
assign Coef[125] = 'h12181AA176625EA511A5046DC22361;
assign Coef[126] = 'h6C9E46B9A0357611377D2088286F36;
assign Coef[127] = 'h0E451AA0A0F7C42212C61A282E698A;
assign Coef[128] = 'h580A5BA02077DC2100C5728837BCB3;
assign Coef[129] = 'h084C05B033EBFCE3B5DF60E840FC0A;
assign Coef[130] = 'hF2FA5FFFDC56DD7A71138CDF01417D;
assign Coef[131] = 'h27FA19E9CC3C3C6E14B69C8F134779;
assign Coef[132] = 'hFFE0437ACC9C31E3E8A53CCF19106C;
assign Coef[133] = 'h3433004B45102BD2909216FF52966D;
assign Coef[134] = 'h3A774513C4841B7B87235CDA44F6DE;
assign Coef[135] = 'h70A31A02A5033AC637933F9D1F8C9E;
assign Coef[136] = 'h6AD11F97A56FDD6B875F0ED9F13A1C;
assign Coef[137] = 'h7B891F9CB3C7A034A7DE0838BEAD98;
assign Coef[138] = 'h5A7CFD9D324FE87967774E5BF4FC17;
assign Coef[139] = 'h583987BDA2F3DEF20ED36C5BFDE796;
assign Coef[140] = 'h3ECD9DBF20DBF3CB0F5F040DB1FD22;
assign Coef[141] = 'h64FD9B3321EE1C61217F56CD5D78BB;
assign Coef[142] = 'h38AA598DC34EF8221DB6594FD9BD11;
assign Coef[143] = 'h572A1C854504ACEB034F0A5F999031;
assign Coef[144] = 'h6DFB55185CA86840252B8B7E8F86C7;
assign Coef[145] = 'h31B95BD574262A23B43B1D4EDB15E5;
assign Coef[146] = 'h67F21BFC47BC6CC1389E4F9EC3C25B;
assign Coef[147] = 'hE14F4540CFA84C423DC168FF774DD4;
assign Coef[148] = 'h079E8F0C4396F89661051A5E2987F1;
assign Coef[149] = 'hBBEED60FC339384037463ADE198708;
assign Coef[150] = 'hC6DD430B64551EA05BE90A6A07AD2A;
assign Coef[151] = 'h4F0A09351077F0E0537C47A8A77E73;
assign Coef[152] = 'h5448DC3122FF9F6273413A6DA37F83;
assign Coef[153] = 'h42D75BA2B237B7228BFB5B0F07692B;
assign Coef[154] = 'h12800D9122EF5C80BBC50B28B67B54;
assign Coef[155] = 'h5AC14B93338BDDD3357A4388E6AD1A;
assign Coef[156] = 'h51E8653E4C34B8E363B60C9E97454C;
assign Coef[157] = 'h6162404ECE50501B90913CEF12C561;
assign Coef[158] = 'h2422507E4FD83843500516AF43D77D;
assign Coef[159] = 'h7A32484BD69C38F34031147E544361;
assign Coef[160] = 'h7AB6520AD704E89AA70F78BB5C1E7D;
assign Coef[161] = 'h72F74093D0ECBEBB3741189BD68E2A;
assign Coef[162] = 'h51C0159F8167CE7B370A4DE11076B3;
assign Coef[163] = 'h4AC88D87A12BE77883CF6D69A92CAF;
assign Coef[164] = 'h1258978FA0CFFE543F535A49D17C9E;
assign Coef[165] = 'h405D52B520FBBCB647534E7973ED9F;
assign Coef[166] = 'h50FD4BB5A26FCADB59202EB98DEE87;
assign Coef[167] = 'h78808B35036B79B85D462E69136B9A;
assign Coef[168] = 'h6E78991CCA2728D84EA4032A7EB6BF;
assign Coef[169] = 'h4D3B0995D886F27807E84B1FBC16EB;
assign Coef[170] = 'h65331E04D68048C829A94EDE0414E4;
assign Coef[171] = 'h7DFB4594CE2420A8048F0EEF1AD37D;
assign Coef[172] = 'h75E80201D5706EE4148B5C5FD316FD;
assign Coef[173] = 'h75F2035F6D3C3122AC971AD61F9754;
assign Coef[174] = 'h5DCB8C8C858FAF392369301BB04489;
assign Coef[175] = 'h575E460C1805F0A2D168789CE9552D;
assign Coef[176] = 'h67975F84C5DF0C631F677A2C2B25F8;
assign Coef[177] = 'h07CB908D4AABB8C2BCE3181D2276C9;
assign Coef[178] = 'h59CA4F922B23ACA2F9C841796E7802;
assign Coef[179] = 'h1DC1118E93237A022FDA61A8212ECA;
assign Coef[180] = 'h4DCE501D3C639E2228CA1E08A5EF41;
assign Coef[181] = 'h59C5C981032BEEB21767C4B8E67BA2;
assign Coef[182] = 'h71F8435CCC107A81209D3C8F0A5275;
assign Coef[183] = 'h72A20A5F4EC83A7930947CCF48C070;
assign Coef[184] = 'h74A1524F4FC830A9588A14EF445075;
assign Coef[185] = 'h7435180A5788401B808536FF5AD375;
assign Coef[186] = 'h462B9389C40C8839667F5CCB55D63D;
assign Coef[187] = 'h7253039D83680811A7966ACE18F2AF;
assign Coef[188] = 'h53F9D385916CEAB83DA64C09D4771E;
assign Coef[189] = 'h325D939E81EBF4BB4B671B38A3A49F;
assign Coef[190] = 'h0059D51EB1EFDEE1A7424A29B42D8A;
assign Coef[191] = 'h1849B18F206FEA314F470C09E5789E;
assign Coef[192] = 'h58DD92B723EFE83A68FA7C7850E91B;
assign Coef[193] = 'h78E5D11E104A3071586EBF68C3397C;
assign Coef[194] = 'h7EBBCA0ED5AE4EC84CB23BC95A2C80;
assign Coef[195] = 'h5DB5104DD4866478C87A39DF4585E0;
assign Coef[196] = 'h51F1160D6DA06008043A234FC0446C;
assign Coef[197] = 'h6FAD8004DF2000B97EE326AA0442B5;
assign Coef[198] = 'h656B1015DE0038AB10833FA64A11A9;
assign Coef[199] = 'hE1C741055F8C6EA9A2074C4FDC9525;
assign Coef[200] = 'h599B434B5E27AC0B2C465B3FF81FC0;
assign Coef[201] = 'h3D8DD304B1C50E41932A6EBFE084A3;
assign Coef[202] = 'h7D8D0B01E643C4610F7F4BC9060380;
assign Coef[203] = 'h2FC9129CBE06F6AB60AA588D2F7FF2;
assign Coef[204] = 'h2D9D47903A23C50057444848213726;
assign Coef[205] = 'h55C9139838AAFE0127660B58AF1C43;
assign Coef[206] = 'h1DD352823BAFDE0131E65B09A6BB53;
assign Coef[207] = 'h31C1529291AAA8A17B6C43B8EFADC2;
assign Coef[208] = 'h21AC2154C49C23BB68976D8782107D;
assign Coef[209] = 'h672CD91DDE887895089B7CAF064275;
assign Coef[210] = 'h67A458CD4448288A581B14EF464265;
assign Coef[211] = 'h24335018D6C838BB445B74AF485075;
assign Coef[212] = 'h607D130FD78964D9A6924E8B14D6B4;
assign Coef[213] = 'h5B4BA387C06896AA57224383D6D434;
assign Coef[214] = 'hA1DB9117826FCCD3776A9BE8B0FC9A;
assign Coef[215] = 'h1B59831F03EFCF631F1709E9F0BD1F;
assign Coef[216] = 'hD9493797A06FEF5B2F5346697BAC9A;
assign Coef[217] = 'h4BDCB395B14BED7127C20481E8AD96;
assign Coef[218] = 'h18C993B682EBE8FA51521C29CCE91E;
assign Coef[219] = 'h2DE1D89D826EEAD058526649D078B0;
assign Coef[220] = 'h37FA881DF1A4C8BA4F2E536797A9B8;
assign Coef[221] = 'h1B7710CEDD85065D6EBA532C5E142D;
assign Coef[222] = 'h65BAD2C7DF202A905E2642CFCA876D;
assign Coef[223] = 'h35224807C2842A9A4A357F2E1E552C;
assign Coef[224] = 'hE5A908165D04488A5A3154AE1A03E1;
assign Coef[225] = 'h858B8B46CF00212B5A1256CFD325A5;
assign Coef[226] = 'h65CA5B8E8F85F8622B52458BBAD129;
assign Coef[227] = 'h2D5F1904DC2F98706B5352ACBCBC3E;
assign Coef[228] = 'h15DC538ECA6BA4CB687E70CC68D168;
assign Coef[229] = 'h5F4143015FAFF082597003286EAAFA;
assign Coef[230] = 'h794813138A23C22271E51129EAEF82;
assign Coef[231] = 'h4DCD5394992FFEA3696E796CA33E02;
assign Coef[232] = 'h514919900DE7F822FDEB914D8CBA59;
assign Coef[233] = 'h41D55B8B0FABAE22626F53E03EED02;
assign Coef[234] = 'h35BC211EC40C20D94AD9248E0CC825;
assign Coef[235] = 'h6EB81ACC5480786B481974E71C4235;
assign Coef[236] = 'h76A4089CDCC8282D489B346700537D;
assign Coef[237] = 'h6630901D57880AF9441B7657144225;
assign Coef[238] = 'h7A7E208C50C932D0FEA334EE5CD2BD;
assign Coef[239] = 'h437021CFD3040569F3222092D08AAD;
assign Coef[240] = 'hE95A435E83ECC7EA1D1F39A8DA4EBC;
assign Coef[241] = 'h99CDB38683E7EDF9B3DF2979F0FC8F;
assign Coef[242] = 'h035891978363F5603B472949EAEC0F;
assign Coef[243] = 'h1B5D91BF806BDBF87BC726C1EBFC82;
assign Coef[244] = 'h38982BB698EAD268185306E011E992;
assign Coef[245] = 'h7C644A9618EA62A818F707E11EE8AE;
assign Coef[246] = 'h4FF8881D91265A78481922E9D8ACBC;
assign Coef[247] = 'h475680C4DF8042BBCF7C41CED696A8;
assign Coef[248] = 'h1D6A8806CC046ABB4629B2A78A46FC;
assign Coef[249] = 'h26299A15C12108DACE0924671E412C;
assign Coef[250] = 'h2D2CD216D3C4326A5C1837AE8F42ED;
assign Coef[251] = 'h616C93CED780D006ECB33A1F9E84ED;
assign Coef[252] = 'hD5CF630ED24975620F5F78EF773721;
assign Coef[253] = 'h1BC8D105A90F8588EB13784BD6BE21;
assign Coef[254] = 'h3F1F900BCFA7C6D05469386DCEFF89;
assign Coef[255] = 'h1D4F13008F26966169ED7BE9CEA969;
assign Coef[256] = 'h2B451B079C67EAC04D7703288EAEAB;
assign Coef[257] = 'h1D4559158FAEDC095FE49169ABFD73;
assign Coef[258] = 'h195419968F2FDF2169A7F3A9AA0F4B;
assign Coef[259] = 'h4B440B0B0FA387831D476AF44ABF8A;
assign Coef[260] = 'h35ECA314EE0038D9CE9074860E4025;
assign Coef[261] = 'h67B900DD52C0485FDC9D754710D135;
assign Coef[262] = 'h64A0889C57481AAA4C107E0705D2BD;
assign Coef[263] = 'h5EAB409C52C048FF4C59664718C0B5;
assign Coef[264] = 'h62EC339CF0C538FB6E17769756D2BC;
assign Coef[265] = 'hF14B004F908021B57E97528B52B8A5;
assign Coef[266] = 'hC9CFC34E8169CDE0BF13F3A8623FB9;
assign Coef[267] = 'hE14FB117986FCDABAB177389F1EC9F;
assign Coef[268] = 'hD949233E88EFF721DB732C69F0FD8A;
assign Coef[269] = 'h59D8B3B688EBDD6131F707C8B1FD9B;
assign Coef[270] = 'h09DD33B680EACC3858DF4C01D1689E;
assign Coef[271] = 'h6BF19296996A487C581F47490279BC;
assign Coef[272] = 'h197F1A0688665A3DDE3663EDC324AC;
assign Coef[273] = 'h1D7B0284DC8166B8EFB9524D9AD7BC;
assign Coef[274] = 'h4DBE800CD6010219C49BF14E0E44B4;
assign Coef[275] = 'hA77D9095DA60689C0CDD408F8F51A4;
assign Coef[276] = 'h273CC004D500602E48AFC02F0EC8FC;
assign Coef[277] = 'hC56C934EDE806A4B2B1EF08E55476C;
assign Coef[278] = 'hC1CC910DDA84BD594B9B38AF89D6BD;
assign Coef[279] = 'h494D610FC28AF5B84FD351ACDD0CC0;
assign Coef[280] = 'h1D9F1A84DE86C40A4977538C9B3DE9;
assign Coef[281] = 'h13DB9952CF2277A04925E22CC4BBC8;
assign Coef[282] = 'h19D71B018FA6DF495BFF5128DEAF42;
assign Coef[283] = 'h1DCD1B118E26FD10FF6F7B0C8EAFCA;
assign Coef[284] = 'h5FD71A048F26CD087FEF7169CFBF58;
assign Coef[285] = 'h59554B1F8DA2CF69FB77D22888BF0A;
assign Coef[286] = 'h44AA215E780968DD4A9DA50F92DC25;
assign Coef[287] = 'h64A808DD7AC83AF74818352F05D335;
assign Coef[288] = 'h64A868D55B4808BF4808340717C0F5;
assign Coef[289] = 'h46A8009C72483AFA4C0B240656D2B5;
assign Coef[290] = 'h4EA9208DD2496AFE4E0630AE50D537;
assign Coef[291] = 'h8A4F335741C811F3FA166B89D002B1;
assign Coef[292] = 'hC1C973570B6245E1FB177189F30989;
assign Coef[293] = 'hE14B234F0167E5F9BB972989F1FE9B;
assign Coef[294] = 'hC3D073FE886FC7E0D997ABA1F1EC9B;
assign Coef[295] = 'h8958F3FF88E7C7F1D9572D49F1FD9B;
assign Coef[296] = 'h4B60F0B688EAC7B89946A581507E12;
assign Coef[297] = 'h4970BA1699EA22BCD8570780D3799C;
assign Coef[298] = 'h4F3588DEDCA672BCDE3A03E9CFA488;
assign Coef[299] = 'hCF3A4CCCD58562FBCE3E43AAD686B4;
assign Coef[300] = 'h4CAED0C4D40D4298CE2A1B2ECF43B4;
assign Coef[301] = 'h4E289894514522F95C6E13269E66B4;
assign Coef[302] = 'h6E29D085D78862984CBF412796C2FC;
assign Coef[303] = 'h4729A1CFD90C0B4BC81B5B175B56EC;
assign Coef[304] = 'h65D8BF4FCD88DDCF4E1E22BE45C460;
assign Coef[305] = 'hD5D9BB4FF3EECF49EA5BA92DD92D54;
assign Coef[306] = 'h6DC97A4DCF2E420BEEFE3BA984AFCB;
assign Coef[307] = 'hAD571A46CF26C7024FB77984CBEE48;
assign Coef[308] = 'h59541A559D2ED71269E6DBACDE3D48;
assign Coef[309] = 'hC9403B478FA6BF097FBC49ACCB2D4B;
assign Coef[310] = 'hD3D51A579D26BF4A7D7EFBA8822D4B;
assign Coef[311] = 'h5DD51A169D22FF0BF97571E8C33F5A;
assign Coef[312] = 'h65A8A9D478156A695AD63D061AF334;
assign Coef[313] = 'h66A960957AC97A7F4C193D6713D2B4;
assign Coef[314] = 'h64A948957B480AF84CA8376717D2F5;
assign Coef[315] = 'h56A9A088F3C938FE4A0F67475040B4;
assign Coef[316] = 'h06A1619D61C9A2F74E136B6B5191B5;
assign Coef[317] = 'hC3CB33CF9BA811EADA177BC9F094DD;
assign Coef[318] = 'hD3CBB35F9962C56B7B9E79A1F09D99;
assign Coef[319] = 'hC9CDF3DF89EEF5EBB91689E9F0EC91;
assign Coef[320] = 'h814967FE897AFD40D11699E9F1AC0B;
assign Coef[321] = 'hC94DB3FE287BF5ADD1579DE8F17A93;
assign Coef[322] = 'h3961B8BE18FAE33A91564EE953E899;
assign Coef[323] = 'h0965BAD798E26AFCD8FE4FE1CF78D4;
assign Coef[324] = 'h4FA5A8D7B9ED6ABADC7F4BE1CF0F94;
assign Coef[325] = 'h56B38CCDD585E2BCD63F4BA1DF0184;
assign Coef[326] = 'h5EBDB885D78542BF4E3E4B2D4F00B4;
assign Coef[327] = 'h4E39B895D3096ABF4EFF436D87C2B4;
assign Coef[328] = 'h7E299895F34822FF4E38470945D0FC;
assign Coef[329] = 'h17B9A3CDDBC87A5F4C7F79B95CC2F4;
assign Coef[330] = 'h45DCE9DDD98AEB7F5A9BB1F8DC8FF5;
assign Coef[331] = 'h4FDD6B1D09ABFFCB4BF23BA9D9AF44;
assign Coef[332] = 'h5759F847EF22538968F35BADCF2CDB;
assign Coef[333] = 'h5FD188578D267F185FFFFBADFB1D50;
assign Coef[334] = 'h5BD119D78F26D7085F7EF9ADCD2FC0;
assign Coef[335] = 'hFBD59A479D26F7C8FBF7D9ADCB2E41;
assign Coef[336] = 'h9BD56A5E9FAAD70AFDF7D9A88F2F40;
assign Coef[337] = 'h79D54A1E8FA2EF4AF9FEF9E8CB3F42;
assign Coef[338] = 'h54A928FC601D30FF4E9B39071B62B4;
assign Coef[339] = 'h44A5E8957B4938FE40913F479BD0B4;
assign Coef[340] = 'h76A9E8B4734812FC4CB93F4717D0B5;
assign Coef[341] = 'h7425F09473C912FE4C617F6751D0B4;
assign Coef[342] = 'h5E0DA08CF3499EEFE6F36B1A7190BC;
assign Coef[343] = 'h4BC9F1DEBBC877EFF893FBC1D19699;
assign Coef[344] = 'hABC971DE9BD875AB9997FBA8D08ED9;
assign Coef[345] = 'hAB4B77FF8BFAF561B19699F9F1AED9;
assign Coef[346] = 'hA14B677E88F6D5A0B1978DB9F1ACD9;
assign Coef[347] = 'h99D1F5FEB8F2D520B9D68DE9F07C59;
assign Coef[348] = 'h2945E2FE98FA777C90D79DE1D36899;
assign Coef[349] = 'h7B61EADE99FE62BC5CB64FE1C13A1C;
assign Coef[350] = 'h5F35E8DEBFE562BCD67743E1CF0090;
assign Coef[351] = 'h5F3BFCCDF68562FCC63C4BADCD86AC;
assign Coef[352] = 'h4C35A485710552DEC672632BD980AC;
assign Coef[353] = 'h4E293A9573858A7F4EFF6B21DE52AC;
assign Coef[354] = 'h5EADE8857149327C4E3C6B2F5541FC;
assign Coef[355] = 'h47A9EFFCDD8870ED4AB77B0F5586F4;
assign Coef[356] = 'h6D69EDFFF9887B5F58376B9B598364;
assign Coef[357] = 'h5F4DEBF7A88A5D4BC9F77B89DC2C48;
assign Coef[358] = 'h5F5DFAC58F2A63695AF77BA9D923D8;
assign Coef[359] = 'h1D51DA578D2A57005EFF3B8D9F0DD8;
assign Coef[360] = 'h7B55485E9E26F708DBFF6B8DCD0FC0;
assign Coef[361] = 'hF3575A578F267548FFB6D9ADCF0F50;
assign Coef[362] = 'hDBD35A571D22770AD9FEC9ACCF8D58;
assign Coef[363] = 'hDBD50A5F9EA2BD48DB7FDBE49F1F48;
assign Coef[364] = 'h448868B47A5D90644E2A3B073BA0B4;
assign Coef[365] = 'h64A5E8B463493AF6443A3F679BD0B4;
assign Coef[366] = 'h5CA9B8B1734902F44CB96F071AD0F4;
assign Coef[367] = 'h5C258890734992F44C797F435770BC;
assign Coef[368] = 'h5605E199B34DF6FE66B37B7175F0BC;
assign Coef[369] = 'hB74773CE9BC85BE7FAB33BA9F116D9;
assign Coef[370] = 'hCBC371FF9FF87D4B98B7EBA9F19A59;
assign Coef[371] = 'hB14F677E99FAF5439197A9E8F10C59;
assign Coef[372] = 'hA941757E8CF6F56199C68DE9F12C59;
assign Coef[373] = 'hB955677EB8F2D553B1D68DE8E1E859;
assign Coef[374] = 'h31457EFEB8FB23FC90C605E1037A18;
assign Coef[375] = 'h439578FE38F762FE98DF4FE00F7A98;
assign Coef[376] = 'h5F917ECEBDBD42FED67D4BE1CE9098;
assign Coef[377] = 'h5F1764CCB785227ED6794B69FC06B8;
assign Coef[378] = 'h5E3BE48C730512FDC67863377D00FC;
assign Coef[379] = 'h4E31AC85F309A27E4EBE6B200F32FC;
assign Coef[380] = 'h4E1DFA95734D227E4C7B2B21DDD0BC;
assign Coef[381] = 'h4FBDE9EC7B982A5D46726B274D40EC;
assign Coef[382] = 'h5DCDE96CBA88795F4257A19B590A58;
assign Coef[383] = 'h5FD5F96EABA2F95F52DF7BC959B948;
assign Coef[384] = 'h7D5B685F8B22710952FF2B85CC2DD8;
assign Coef[385] = 'h795578468D2637425EB7BBA5CF0E48;
assign Coef[386] = 'hDB517A5E9D26750A57FFCBAD4F0E48;
assign Coef[387] = 'hD1535B478CA65509F7D6B98DCF0E40;
assign Coef[388] = 'hF9D75A4E8F227D0B599E99E58F2B40;
assign Coef[389] = 'h7BD76A5F9EA23D4B59B6F1E5CFBF48;
assign Coef[390] = 'h6E8C2AB4B85D82754AAABF633BF0F4;
assign Coef[391] = 'h64A5A8B0614D4AF44C386B6399D0B4;
assign Coef[392] = 'h7CB9A8B1614902F44C3137671ED2FC;
assign Coef[393] = 'h4C21B8B163CD82F442617B6158F0BC;
assign Coef[394] = 'h4E85F08DB1CD9A3443F97B6151D29C;
assign Coef[395] = 'hE38760EEBB9C25EFD8B779E37114D9;
assign Coef[396] = 'hA3C3277F9FFC754F98B6DD89E39A59;
assign Coef[397] = 'hA141757E8EF07D6799A68D80E19C59;
assign Coef[398] = 'hE951777E8CF2754799868DA1E15E59;
assign Coef[399] = 'hA951777EBCB27D6591D68DE8237859;
assign Coef[400] = 'h3B55767EBFFB637E90C644A1037A08;
assign Coef[401] = 'h6B353C923DFD6AFE90FE4761085A98;
assign Coef[402] = 'h4B35BECD3FB562FE967E43E10D1298;
assign Coef[403] = 'h0F9334CDB795427EC6794368AD9588;
assign Coef[404] = 'h1E33B484F59DC2F64638632F3D82BC;
assign Coef[405] = 'h4E1DFC84F31D827E4EA863692FA2F8;
assign Coef[406] = 'h5EBDBCA5F15DDAFE46E9632C0D70FC;
assign Coef[407] = 'h4FBCE8EFB99D7A5F443B2B2F5D91E8;
assign Coef[408] = 'h75ECE8EE3899695F40732FEF59A160;
assign Coef[409] = 'h5F5D3A6EBFA6794F42D6ABA54DAB40;
assign Coef[410] = 'h7FD5786B8EA6735EDAD72B854D1848;
assign Coef[411] = 'h7F551A4B8F2635C156FE83858E0D48;
assign Coef[412] = 'hF9575A4F9D267559DFF7C9AC8F0A48;
assign Coef[413] = 'hDBD75A4E8E267D5BDB9EE9ED8F0E40;
assign Coef[414] = 'hDBD47A5F8E223D4ADDDEA1AD0F0E40;
assign Coef[415] = 'hFBD66A4E9FA2BDCBD49EE1E58F1F48;
assign Coef[416] = 'hC48868B5391D82744AB02B23BBE0D4;
assign Coef[417] = 'h64ADE8B1635D9A744C383B63BBF3FC;
assign Coef[418] = 'h7CB9B8B1615D82B44AB91F65BFF0FC;
assign Coef[419] = 'h5C11F8B121CC82B446792F615CF19C;
assign Coef[420] = 'h4685FABD33CDCA7E62317B6158D6D8;
assign Coef[421] = 'hEB8DF2EF1BDC72EE90B3FB2BD192D9;
assign Coef[422] = 'hA345666E9FDC6D4F9886FDA301D259;
assign Coef[423] = 'hA3C3657E9EF87D43B1868DE1A11C49;
assign Coef[424] = 'hA1C3777E1EF2754791868DA121C851;
assign Coef[425] = 'hABC5777E9EFB7DC791C68DE0826B51;
assign Coef[426] = 'h2945F43E3EF3457E90C694E00B7A19;
assign Coef[427] = 'h7B35B4BA37FD0AFE9CCC07600E5098;
assign Coef[428] = 'h1FB7748DBD958AFE967D43612C1308;
assign Coef[429] = 'h5F17B4C9B59DE2FF86796323AC9688;
assign Coef[430] = 'h4C913C80F59DF2F626282B2F7D00B8;
assign Coef[431] = 'h5E14FE91371D827E46E9636C2DB2C8;
assign Coef[432] = 'h5E39B8A5E31D92F406F9EB250DE0D8;
assign Coef[433] = 'h7EBCB8EDF39D427F460127275DA2F8;
assign Coef[434] = 'h5A9CE86F2898787750432FCF4DB340;
assign Coef[435] = 'h74DDF86DB4AF7D6748C7ABE31CA040;
assign Coef[436] = 'h7FF3384E8EA45345C0AEABEF0F0048;
assign Coef[437] = 'hFB577A438E244251D2DEAB8F0C0948;
assign Coef[438] = 'hFBD75A4E9DA6BD4BDFDE898C0E0C48;
assign Coef[439] = 'hBBD77C4F9E267D4BDF96A9AF0F0F41;
assign Coef[440] = 'hF9F37A4F1E263DCFD89EF98D0E0B40;
assign Coef[441] = 'hFBD65A5F9EA22C4BF89CF1A40E1F40;
assign Coef[442] = 'hE498FEF4295D826C6AA82B03BB70D0;
assign Coef[443] = 'h4CB9FAB0215D82744A310B69F9F1FC;
assign Coef[444] = 'h5C39B8B0615C82B448F95F655EF1FC;
assign Coef[445] = 'h5C15F8B1A1CDC2B040715B61FDF3D8;
assign Coef[446] = 'h4E85F8B9B3CD4A7C627B7B69DDF3D9;
assign Coef[447] = 'h638170EFBB9C2B6F98B1FFEBF9D659;
assign Coef[448] = 'hE3C7766E9FF82D6F9094FDEB03D359;
assign Coef[449] = 'hE1C3756E9EF86D4FB984ADAA81DA59;
assign Coef[450] = 'hA346777E9EF07D479986ACE2AB1A41;
assign Coef[451] = 'hE347777EBEB36D4791C6ACA2031A49;
assign Coef[452] = 'h6B45763EBEF3286E90C6CCE00A7A09;
assign Coef[453] = 'h6A35F6933FF5027E94EC45600E5219;
assign Coef[454] = 'h4A97B681B7D5EAFEB66C42202E1389;
assign Coef[455] = 'hDE96B489B795CAFFA730EB26AC9688;
assign Coef[456] = 'h5E11E480B51D82F4266923362C50A8;
assign Coef[457] = 'h7E1DB4B0379DA27406E96B682EB288;
assign Coef[458] = 'h5E3CB6A1A75D82FC06E96F216D70C8;
assign Coef[459] = 'h5CB4B8A922DD2A7504616F0F0CB140;
assign Coef[460] = 'h5EB0F8E82A9D2C674047AF474CB140;
assign Coef[461] = 'h53D57A7CBE97617750C5EA870DB140;
assign Coef[462] = 'hDF773C4F9C8501CED4C7AA870F0240;
assign Coef[463] = 'hDB773E4ACCB420409686A9070E0440;
assign Coef[464] = 'hFB577E4F9FA6345AFF9FE98E0E0E40;
assign Coef[465] = 'hFBDA7E4F9E253D4FFF9CA98E0E0740;
assign Coef[466] = 'hFBD67A4F9EA47DCFFC9CF88F0F0B40;
assign Coef[467] = 'hEBF61A4F1EA22CCFB48DF0870F1F40;
assign Coef[468] = 'hE09BEEB0A317926020AA0F2B3A61D0;
assign Coef[469] = 'h6C31B8B021DD923448315B61F9F9DC;
assign Coef[470] = 'h7E39B8B0615CC2304A7B5F617DF1FC;
assign Coef[471] = 'h5C1598B021CE823442715B615CF1D8;
assign Coef[472] = 'h5A15F0B831CCD67CE2717B6179F3D8;
assign Coef[473] = 'h23B5F0EFBF9C0A76C031FD6F491359;
assign Coef[474] = 'hA3C1746F9FD86D4F1884FDE383D779;
assign Coef[475] = 'hA1E7777E9ED03D479086EDABA9D249;
assign Coef[476] = 'hE1E7677E9EB07D4F9886ADE283DA41;
assign Coef[477] = 'hA1E7777EBEF33D4F91C68CA2035A41;
assign Coef[478] = 'h23C5763B3AF3245E90CE4CE0027A09;
assign Coef[479] = 'h7A25B6317E71827E94EE44602A5299;
assign Coef[480] = 'h4A95B481B755CEFCB7784820AC1209;
assign Coef[481] = 'hD29EE408B795EAFFA7796B2AADB689;
assign Coef[482] = 'h5E94B480A79582F52679232FFDB098;
assign Coef[483] = 'h5E11F6A1359DE6F427E96B092DA28A;
assign Coef[484] = 'h5C9DB4B125DD827407E16F692C7098;
assign Coef[485] = 'h5E94F8B8269522F540432F270DB0C0;
assign Coef[486] = 'h70AC787A2291687E0041AFA62DB140;
assign Coef[487] = 'h5AF57C6916B72877D247AEA70C3B40;
assign Coef[488] = 'hFFF73C4ADE9544D1D2CF2EA70F0160;
assign Coef[489] = 'hFB735E4A5CB47DD190DFAA8E0D0040;
assign Coef[490] = 'hFB577E4E9EA575D3BF9EE88F0F0F40;
assign Coef[491] = 'hFBD73E4FDEB43DCBFF9EA98E0F0761;
assign Coef[492] = 'hFBF67A5F9E243C4FFCDC688E0F1341;
assign Coef[493] = 'hFFD77A1F9EA02CDEB49CE8C60F1B41;
assign Coef[494] = 'hE8973EB5915E8724E9AA9B23BB6DD8;
assign Coef[495] = 'h5C3DBEB0215FD23462335B61BDE9D8;
assign Coef[496] = 'h5C11B8B1A55F82B040F95F61FEE1D8;
assign Coef[497] = 'h5C15B0B021EF82B040715B61FDF9D8;
assign Coef[498] = 'h5A15F0A9A19D0E34C2715B6159F358;
assign Coef[499] = 'hEAB574EF3F9C286E9031DDE789D779;
assign Coef[500] = 'hE3A5766FFFD8356F10BEFDEF815379;
assign Coef[501] = 'hE1E7656FFED07D4F9084FDAEA3D369;
assign Coef[502] = 'hE3E6777F1E307D4F9886BDEA83DA61;
assign Coef[503] = 'hE3C5667FFE712D4F98CEACE2235A43;
assign Coef[504] = 'h23457633BA732C4E90CECCE0027A09;
assign Coef[505] = 'h6A25B6317375C2EE14DC46602A72B9;
assign Coef[506] = 'h5AB7B681F755CEFEA6696068AC9289;
assign Coef[507] = 'hDA9FF401B795C6FDA7716A2AECB699;
assign Coef[508] = 'h5C14F481355DC2F027716325753188;
assign Coef[509] = 'h5A1596B025DFE6B407694A692D628A;
assign Coef[510] = 'h5E1DF6A0255FC2B426F946692D2198;
assign Coef[511] = 'h7EBCF8B867DDCA7404432F672DB200;
assign Coef[512] = 'h52B4AA283293A87650412E6F09B140;
assign Coef[513] = 'h7285786A36B3A9F732C62E230DB040;
assign Coef[514] = 'hDAB76C4ED6B465CF8EC6B88F0D1161;
assign Coef[515] = 'hFBD7F64AC61575D892DEA88E0B0342;
assign Coef[516] = 'hFBD77C4FDE357CDBB2DE788E0F1362;
assign Coef[517] = 'hFBE77E4FDE253C4BFF9CF8CE8F1261;
assign Coef[518] = 'hFBE77E477E202CCF9C9CF8C70F1A61;
assign Coef[519] = 'hFBE77A4FD6202CDFB8DCF88E0F1361;
assign Coef[520] = 'hC83F1EB4259D8734E1AA8F21A96998;
assign Coef[521] = 'h5C39BEB0C55EC23061735F61ADE9D8;
assign Coef[522] = 'h5E3994B0457E82B044735F61FEE9D8;
assign Coef[523] = 'h581598B825CEC2B440715B615C6998;
assign Coef[524] = 'h5A15FABD25D66734E0735B6159F158;
assign Coef[525] = 'h6AA772EFDFDC281F88037D6F0DD3F9;
assign Coef[526] = 'hE3AD677FFE5C3C4F380EFD2F09D369;
assign Coef[527] = 'hE3EF677FFED03D4F1084BCEE8B5361;
assign Coef[528] = 'hE3E7677F7EB02D4F980EBD86835261;
assign Coef[529] = 'hE3E6637FFAB12D4F98CE3CA2035A67;
assign Coef[530] = 'h62E57633B273284E1CCE4CE0037A0F;
assign Coef[531] = 'h62013631F3758AEA1CCC4C60A2728D;
assign Coef[532] = 'hDA9FB701F755CAEF37684868AC3389;
assign Coef[533] = 'hDA9F7541B715EEBFA7716A38EDB619;
assign Coef[534] = 'hDA1EF420A59D82A427710A3974A488;
assign Coef[535] = 'h5A1DF6312757E7A4266152282C2B0A;
assign Coef[536] = 'h5A15B6B0A55FC6B427F36E682CB99A;
assign Coef[537] = 'h5CB4EC2C64DFAAF404702F6F2DB001;
assign Coef[538] = 'h50A4682D769B287400512E2B09B303;
assign Coef[539] = 'h76A56E6F76B3EC5F34C72CAA0DBA03;
assign Coef[540] = 'h17E7744ED61579DF87D4788E0D1363;
assign Coef[541] = 'h7FEF664CD63539CFD7D4388E291362;
assign Coef[542] = 'hF3EF4E47FE35FCDFBFDE688E8F1661;
assign Coef[543] = 'hE3EF464FFE157C4BFF9C788EAF1721;
assign Coef[544] = 'hE7E76647FE352CCFFCDC788F0F1321;
assign Coef[545] = 'hE7E76A07F6212CCEBC9C78CE0B1301;
assign Coef[546] = 'hC03FBFB445BF8730A46AC3232D6DB8;
assign Coef[547] = 'h5831B4B045FF82B060735B65AC69D8;
assign Coef[548] = 'h5C39BCB045FE82B005F35761BC68D8;
assign Coef[549] = 'h58159AB825EF82B081735361CD7998;
assign Coef[550] = 'h5A15F0BF25FA2AB4A0535A6149B918;
assign Coef[551] = 'h66B57AED7F98282E0008FD6FA8D379;
assign Coef[552] = 'h67AD676FFE5D784F08087C2729D37D;
assign Coef[553] = 'hE3EF657F7E50394F188CBD8F83D365;
assign Coef[554] = 'hE3E6657F7E903D4F188EBC8E035367;
assign Coef[555] = 'hE3E6665FFA212D4F188EAC8E035A67;
assign Coef[556] = 'h62E564113A6BAC4B18CE5CC0A3FAAF;
assign Coef[557] = 'h620DB7B1FB7DA28A37CA5C002272BF;
assign Coef[558] = 'hB29FA701B755CE9C27585818A8B7AF;
assign Coef[559] = 'hDA9FF545B51DCEBD27516A39F9B51B;
assign Coef[560] = 'hD817D52C251FC3B427614B3875B58B;
assign Coef[561] = 'h9A3FB5A125DFABB023CBDA79252B0A;
assign Coef[562] = 'h5A19B43125F7C2B027E34E69AD3C0A;
assign Coef[563] = 'h5CBD7CA964FFAAB004410F6B21B123;
assign Coef[564] = 'h70A5460D36E3AC7E09423E6BA9BB03;
assign Coef[565] = 'h62A5464836F3ACAE28865C4B0D1327;
assign Coef[566] = 'h17EF444DD681B8DE87D47C4E091225;
assign Coef[567] = 'hE7E3440ED6253CDEE698788E081267;
assign Coef[568] = 'hF7AF6445FE1520CFD79CF8CEAC1625;
assign Coef[569] = 'hE3EB664FDE152CCFDE9E788F0F1665;
assign Coef[570] = 'hE7E76E45FE203C4FDC9C788E0B1325;
assign Coef[571] = 'h26E76A45FE202CDE3C9C78C68B1321;
assign Coef[572] = 'hD1B61FB76DDF9730FF4AD36D2F2998;
assign Coef[573] = 'h1833BEB245FFC3B0E97B9761ACE9F8;
assign Coef[574] = 'h5E119CB0C5FFC2B025FB57612468DA;
assign Coef[575] = 'h5A119AB805EB82B080E3526105F85A;
assign Coef[576] = 'h5AD5F8BE258AC59C404BD8ED01B919;
assign Coef[577] = 'h67AD68ED7E99285E40087D6F89F379;
assign Coef[578] = 'h67AD67FDFA18284F2E48FD6F2BD37F;
assign Coef[579] = 'hE7AE677F7A102D4F388CBD8E8BD367;
assign Coef[580] = 'h67AE677F7A18284F188EBC8E83D367;
assign Coef[581] = 'h63E64757FA212C4F188EB48E22D327;
assign Coef[582] = 'h63856651FA63AC4E1DCED448A27AAF;
assign Coef[583] = 'h620F9691F3558A0C2FCA5420A263BF;
assign Coef[584] = 'hD29FB701B355C68D277A5878ECB78F;
assign Coef[585] = 'hDADFB54DA715EEB52751F279F5B51B;
assign Coef[586] = 'h5A1FB4202555C7B42753DB797DB59A;
assign Coef[587] = 'hD217B7310577C7B023C3D169A1A90B;
assign Coef[588] = 'h581D9531A5FFC7B007E34E682D3C0B;
assign Coef[589] = 'h5EBDD4A467FB8AB003430F69219947;
assign Coef[590] = 'h50A5E42936E3E8A501424D6A013303;
assign Coef[591] = 'h7EA7664972E928F610845D6B09BB07;
assign Coef[592] = 'h76AF6645D6212C4FA7C25C9E019325;
assign Coef[593] = 'hE7AFCC47D6057CDFE3CE781E111727;
assign Coef[594] = 'hE7AB6645DE05ACDFDF8C799F2B0625;
assign Coef[595] = 'hE7EF2F45DE157CCFFE98799E8D1625;
assign Coef[596] = 'hE6AF6E45FA14ACCEFE9C79CF8B1325;
assign Coef[597] = 'h66AF6E057B012CDEBE9C784F8B9325;
assign Coef[598] = 'hD8139EDE4D898714FCCAD5EDA74D38;
assign Coef[599] = 'h1E339CB0C5FFC3B0E4F3CF61AC68BA;
assign Coef[600] = 'h1A1196B045FFD3B085F35F61A46859;
assign Coef[601] = 'h5C1590BA45EBC3B045F3D261297858;
assign Coef[602] = 'h5AD5FA7E34AB30BC445259ED2DB959;
assign Coef[603] = 'h66A568FD7E99781C041A7D6F2DB1B7;
assign Coef[604] = 'h67AF67F5FA19384F2E0AFD4FAEF3F7;
assign Coef[605] = 'h67AF6F757A183C4F080CBD0E8BD367;
assign Coef[606] = 'h67AE6F7F7A38294F180EBC868BD3E7;
assign Coef[607] = 'h67A667557A212C4F380E348EAA73A7;
assign Coef[608] = 'h630746D1BB6BAC4E1D8E744CA2FBBF;
assign Coef[609] = 'h630F3711B37F86CC2FEA5044A263BF;
assign Coef[610] = 'hFA1F9741A155C688277BF038F5B79F;
assign Coef[611] = 'hDB1FD74D2515C7942753F179F4B58B;
assign Coef[612] = 'hD817B56905D6C7902753D379F5B51B;
assign Coef[613] = 'hFB55D733857BC7B427C3D56825B90A;
assign Coef[614] = 'h1A579730847FD7B027C3D76921391B;
assign Coef[615] = 'h5C1DF7A0647BEAB00142076929B927;
assign Coef[616] = 'h60E6FE50266AA8BE23C2186B21BB27;
assign Coef[617] = 'h40AFEE206661E8BD0BC65D6A09BB27;
assign Coef[618] = 'h66EFE544C20178FC93825D3E919327;
assign Coef[619] = 'hE7AF4741DA1534D9878A78DE719227;
assign Coef[620] = 'hE7EF6745DA1D7CCFEF8C799E5D8727;
assign Coef[621] = 'hE7AB6E45DA157CCFFF98F99EF99725;
assign Coef[622] = 'hE6AFEE45FA153CCAFA9879CF0B9325;
assign Coef[623] = 'hE6A76E015B012E4E7E9C594E8B9325;
assign Coef[624] = 'h9C339EDEED9F97B8ECCA9D65AD4936;
assign Coef[625] = 'h18519DBAC5B3D3B0C6D2D96DA86819;
assign Coef[626] = 'h1A1194B2C5F357B08DF35F618C685A;
assign Coef[627] = 'h1A559ABE24A353B0C4D3D1E1257819;
assign Coef[628] = 'h5AF538FE64A3509C7052D9E581F933;
assign Coef[629] = 'h74A5CAFD7B19F87C4C5A7D6FADF1F7;
assign Coef[630] = 'h64AFEFF57A59BC4F6C0A754FADF3F7;
assign Coef[631] = 'h65AF4D757A10384F280ABC1F8FD3E7;
assign Coef[632] = 'h65AA4F757A18384F180EB50F8FD3E7;
assign Coef[633] = 'h67A663D5FA28384F3C0E340E8FF3E7;
assign Coef[634] = 'hE6074711BB238C4A398ED04CA67BAF;
assign Coef[635] = 'hF30B97B13377C4082FEAD144A66BEF;
assign Coef[636] = 'h8B1FD741A117D79D275BD059FDB59B;
assign Coef[637] = 'hCBDF954FA115F7B56753F179F5B59B;
assign Coef[638] = 'hD857956E05DED3902353D168F19D1B;
assign Coef[639] = 'h5B579532857BC79027C3D578C0391B;
assign Coef[640] = 'h9855B532247BD7B023D3C769292D1B;
assign Coef[641] = 'h5835F724447B86B023D20768A9B997;
assign Coef[642] = 'h6CA5E6A07F683E3C02961D6D89BB27;
assign Coef[643] = 'h64AFCFC0E27BADFC3BC6DD6A81BBA7;
assign Coef[644] = 'h4EAB5D45C215FCFA8B82537E9997A7;
assign Coef[645] = 'h6FAB6745D07D36DEF38A791E591727;
assign Coef[646] = 'hE7ABC745FB1D3CCBEF98F99ED99324;
assign Coef[647] = 'hE7AF6F47BB1DFCCFEF98B91FD99725;
assign Coef[648] = 'h67AFE641BB7C2C4F7E9E79CFBF9325;
assign Coef[649] = 'h66A72E05FB412ECE7EB8794E9B93AD;
assign Coef[650] = 'h9F311F5EEC9995B4F5C299EDAF3835;
assign Coef[651] = 'h1811D4BAC4E3D790DDD2DDEDAF4819;
assign Coef[652] = 'h1A5196B6C4F3529085F3DF6188285B;
assign Coef[653] = 'h1A55D8BEA4AB52B091D7D0E181381B;
assign Coef[654] = 'h5EF5D87EF4ABF89C5056DDEF81B971;
assign Coef[655] = 'h64B5EDF5EA19585C6C1A5D6F8DF1F7;
assign Coef[656] = 'h65A7CFF5FB59384D6E0AB54FAFF9F7;
assign Coef[657] = 'h65AE6BF57A18384F680A3C1F87F3E7;
assign Coef[658] = 'h64AE4BF57A18384F2C0EB40F8FD3E7;
assign Coef[659] = 'h66A66BD17B28BC4F2C0EB006A673E6;
assign Coef[660] = 'hE60703D1BB2E9C4E3DAED04CAF6BFF;
assign Coef[661] = 'hF31F97F1A13C95082F8AD74CA64BBF;
assign Coef[662] = 'hCB5FF741A11FD599275BD05DFCA51A;
assign Coef[663] = 'hD85FB54F8097D5916753D15DF5B51B;
assign Coef[664] = 'hD856B56E04B2D1B4A7D3D3F5F1BD1B;
assign Coef[665] = 'hDA579726A57AA79003C3D4E9A1B91B;
assign Coef[666] = 'h185BB5336473D7B093D7CDE170AC1B;
assign Coef[667] = 'h5899D5A02579D2B043E28778B1B9F7;
assign Coef[668] = 'h4CA7EDA10D783CB830964569819BB7;
assign Coef[669] = 'h646FEFA0CB78BCFA5F8ED56D81BBA7;
assign Coef[670] = 'h642BDDC5E30874F8C396D17ED987A7;
assign Coef[671] = 'h620BA785FB5D72C9E3AA3D1E5983A5;
assign Coef[672] = 'h67AF2F47FB55345BE398B95FD58734;
assign Coef[673] = 'hE3AB6747FB1C7C4FEF98B99EF99725;
assign Coef[674] = 'hE6AF6F45FB5C3C4E7E98790DDF83B5;
assign Coef[675] = 'h66A7AEC1FB582E6A6AB8714FBF93BC;
assign Coef[676] = 'h55115D5EECB1B59CDFDE194FAF5C33;
assign Coef[677] = 'h1E55D51AE4EB1590D7D6D569AC6C17;
assign Coef[678] = 'h1A11D23AA4E3569091D3DF6D88481B;
assign Coef[679] = 'h1A51D23EE4A3D190D1D659E9883813;
assign Coef[680] = 'h1ED5F8FDBABBF8DC50D6D8ED89B153;
assign Coef[681] = 'h6CB5EBF56A39F87C6D1AB36FADF1F7;
assign Coef[682] = 'h64AD6FF5EB59B85C6E3AB75FAFF1F7;
assign Coef[683] = 'h65AC6DF5FA18B84F6C08B51F8FF1E7;
assign Coef[684] = 'h64AC6BF57B18384F6C0A351F8FF3E7;
assign Coef[685] = 'h64AA4BD1FB2ABC4B2D2AB01FA773E6;
assign Coef[686] = 'hE74F03D19B3E9D4A3FAEF21CAE6FDA;
assign Coef[687] = 'hEB4F97718937D5492FDAF24CF66DFA;
assign Coef[688] = 'hDB5FB7438117F5D96753F15DFCBD1A;
assign Coef[689] = 'hD9DEF54EA095F59D675399FDF9BD1A;
assign Coef[690] = 'h9857F76E09923194E75391FDF19D19;
assign Coef[691] = 'hDA57D777897AF59897D790E981291B;
assign Coef[692] = 'h9A5FD5228073D5B0B3D68CF9592C1B;
assign Coef[693] = 'h1C55D5A10C7B56B013F6857D91D953;
assign Coef[694] = 'h6267DFA3E178B9B8B1B6D279819BB3;
assign Coef[695] = 'h6203EFA1F37BB2DB3386DD6899BBB3;
assign Coef[696] = 'h6A2B4FE191593DFCE3BA105E5993A5;
assign Coef[697] = 'h66EBCF879B59F0DDE38A1A9E5987A4;
assign Coef[698] = 'h61ABCF43BB5DB44BE71E3B1FDD83A4;
assign Coef[699] = 'hE6AB67C7BB5DFC4FE798B99FFD87B4;
assign Coef[700] = 'h66AFEFA7BB5C3E6EE2BC7B0DDB83BC;
assign Coef[701] = 'h66A7EE83FB5D2E6EF6B9731DFD97BC;
assign Coef[702] = 'hC1495E5CB803B5D8F79658CFA93D71;
assign Coef[703] = 'h1E51D77CECA355D0DEDE5D6DA90813;
assign Coef[704] = 'h1E51D638A4E350909FD75FE98A4853;
assign Coef[705] = 'h1A51F23EA4235198D1D6D9E98B3813;
assign Coef[706] = 'h1EB5EA77B82BD8DC59D2D96DABB953;
assign Coef[707] = 'h64B5EBF5E839F85C6E3A3B4DA9F9F7;
assign Coef[708] = 'h64A9CDB5E91DB05C6E1A3F5DBCF1F7;
assign Coef[709] = 'h64AA6DF56B18B84F6C0ABF1FAFF1F6;
assign Coef[710] = 'h64AA4BF55B38384F6C2AB70FAFF3E6;
assign Coef[711] = 'h64E24BD55B3ABC4B2D2EB21FAEFBE6;
assign Coef[712] = 'hE7474BD39B3E954B3F8EF21DBE6BCA;
assign Coef[713] = 'hE34F1773893E9549279AF04D7649DA;
assign Coef[714] = 'hDB5EC56B881FD515EF53F9D9FDAD1A;
assign Coef[715] = 'hD9DFF54E809FF5D5E753B9F9FDBD11;
assign Coef[716] = 'h9856FD6A08B27190E7D7D1F9799C13;
assign Coef[717] = 'hC857F76BE8FA319997D7DCF9153919;
assign Coef[718] = 'h0B55D76E8473159893D6C8F9702C53;
assign Coef[719] = 'h5E3BFDA66D7A11B083F68769D95877;
assign Coef[720] = 'h6829DDA3C972BCB8A3F6C77D999FB9;
assign Coef[721] = 'h622FEFA39B79BBF5B3B6DC7D99F1FD;
assign Coef[722] = 'h222BDFE7C358F0F8E332FEF8D99DB4;
assign Coef[723] = 'h4E2FEF87B95971FDE3BAFD1C79A7B4;
assign Coef[724] = 'h626F4F67AB5D7469E738FF1DFD87B4;
assign Coef[725] = 'hE6ABEFC7FB5CFE6FE618BB9F7997B4;
assign Coef[726] = 'h668FEE87FB5C166AE2B87F0D5D87FC;
assign Coef[727] = 'h66A7EFC5D359B66EE6B9731DFD97BC;
assign Coef[728] = 'hC04BC1DCB80F35DCEF3295EFAF5411;
assign Coef[729] = 'h1D51D110E02314909BD4DBED8A2813;
assign Coef[730] = 'h1E53D23EA4A351909BF75DCD820853;
assign Coef[731] = 'h1A55501FB423509CD1D6D9C58B1813;
assign Coef[732] = 'h5E91F275F82B70DC43D6D94DAABB73;
assign Coef[733] = 'h6CB9EFB5E83BD87C6E32BB6FADB9F7;
assign Coef[734] = 'h642BCDB5E97B90746F3AB75DBFF1F6;
assign Coef[735] = 'h64AA6FF5EB18B86C6C2ABF1FBFF1E6;
assign Coef[736] = 'h64AC6BF5DB3A984D6C2AB21F3FF3E6;
assign Coef[737] = 'h642A4BF5DB3A994B6D2EB21FBEEBEA;
assign Coef[738] = 'hE74A4BF3C93E95493DAEF385AE4BCA;
assign Coef[739] = 'hF74F4F33C93E95492FEFF21DF64DEA;
assign Coef[740] = 'hD35ECF6B889FF5596753E9D97DAD13;
assign Coef[741] = 'hD95E7D4EA89FF5D1E753B9F9F9BD10;
assign Coef[742] = 'h5874516E88B8119057D3DDDD799D53;
assign Coef[743] = 'h5A53C76B89FA35D895D7DCC93C0859;
assign Coef[744] = 'hCB57D77A803A35D1B3D6DCE9718C53;
assign Coef[745] = 'h5859DCB2E57911B093F68F5999CC55;
assign Coef[746] = 'h4837DEA22178ACF1B3FEC469DBF1FF;
assign Coef[747] = 'h666DCFA3B378B1F9B73EC6F9F9B3FF;
assign Coef[748] = 'h42294DE7B158BFF9E330DF7979C1BC;
assign Coef[749] = 'h660BCFE2B959F67DE630FF39F9C5F4;
assign Coef[750] = 'h672BEFE7E15CE269E732FF397DE5BC;
assign Coef[751] = 'hE5AB6FE7FB5CFC6DE73AFF3F7DE5FC;
assign Coef[752] = 'h66AFAFA5FB5C1668E6B8FF09FD47BC;
assign Coef[753] = 'h66A7EEC1EB599628E6B9F739FDD7FC;
assign Coef[754] = 'hD041424CA82315DEC39E99CF8F5871;
assign Coef[755] = 'h1E51D214B42355D4DBDAD9CF894813;
assign Coef[756] = 'h1F51D216A42116D0D3F75DCD8A0857;
assign Coef[757] = 'h1A55F255B42314DA53D659CD8B1853;
assign Coef[758] = 'h54956275BA32B8DE5AD6DDCF8BBB53;
assign Coef[759] = 'h54B5EFB4E03B927C6F3ABB5DAFF9F3;
assign Coef[760] = 'h742A4FB1E47B907867222F1DBFE9F6;
assign Coef[761] = 'h64AE4FF54D38BA6C6C2ABF1FBDE9F6;
assign Coef[762] = 'h64AA6BF54D5E8A6C6C2AB60FBFF1E6;
assign Coef[763] = 'h666E4BB54D3A81496C2EBA1D2ECBE6;
assign Coef[764] = 'h676E4B33C93C95493DAEE2952E43CA;
assign Coef[765] = 'hE36E4B73C9389549A7CFB29D7C4DD2;
assign Coef[766] = 'hD35E4F6FA0BBF55967D7B9D97CAD12;
assign Coef[767] = 'hD0DE4D4EA8B375D1E757B9DFF99D10;
assign Coef[768] = 'hD0747D6A88B971D0D7D58DEB518951;
assign Coef[769] = 'hC2757B7AF0FA35D8D0D6DCC95B0953;
assign Coef[770] = 'h8351736BA8BB35D1B1D6CCC9582C13;
assign Coef[771] = 'hD259DBB3A47A1598D1F6C5E99B695B;
assign Coef[772] = 'h6E7FDFA3B578B5F9D0BECCEDF3F5FA;
assign Coef[773] = 'h421D4FA3E168B5F9F23ECCBDDBE7FF;
assign Coef[774] = 'h626F5BE7B9C8B9EDE335DE39F9D7BC;
assign Coef[775] = 'h632BCBE3A9D96578E732FE19FD45DC;
assign Coef[776] = 'h6A2BCFE389DCC568E631FF397DF7DE;
assign Coef[777] = 'hE3AF6FEFB9DCF569E730FF3BFDD7BC;
assign Coef[778] = 'h672FEFE7E95CD668E6B17F1D75C39C;
assign Coef[779] = 'h6E27CEA38959B668E6B15F3DFDD7FC;
assign Coef[780] = 'hC00943D4B80795DACB909BCFDD4C51;
assign Coef[781] = 'h56115355B42754D2DBDA5FDB8A4817;
assign Coef[782] = 'h1B535217F4611590D3D75DCF8A0853;
assign Coef[783] = 'h52577257B42035DA53DED9CB8B0A53;
assign Coef[784] = 'h56F56255FE2239DE4A9EDFCDABBB73;
assign Coef[785] = 'h5CB24FB5EC7B92786F32AB5D3FF976;
assign Coef[786] = 'h5CBA6FA5E47B93706C32AB1D3DE9D6;
assign Coef[787] = 'h64AAEDA5C5389A606E2AAB1DBDF9E6;
assign Coef[788] = 'h64A84FB54D7A9A6C6C2AA71D2FC1E6;
assign Coef[789] = 'h642A4BB35D3887496D2EA31D2E49E2;
assign Coef[790] = 'hE76E4B93C93C9549BDAEBB1D2ECFEE;
assign Coef[791] = 'hD6624BA3CD381549FFCEE08F744942;
assign Coef[792] = 'hD9566D6F8099B559F7C7A19B7C8D12;
assign Coef[793] = 'hD0D64D6E0899F5D5F35499DB799C11;
assign Coef[794] = 'h5074546A88B039DCD2D7CCCB598C51;
assign Coef[795] = 'h62477B7ED0FA15D8D1D7FCCB114A51;
assign Coef[796] = 'hC353522FB8F235D9F1D68CD9590C51;
assign Coef[797] = 'h5B51DEA2E47297D091FFCCC9E94057;
assign Coef[798] = 'h4A77DFA3F56814F8F0BECD3BF9EDD8;
assign Coef[799] = 'hE26B4AA3A16A97F8F13AC629BDFF9A;
assign Coef[800] = 'hE26948EFA1DA8568E731CF3A79E598;
assign Coef[801] = 'h67496FEFB9DFF768C131DF2BFDE55C;
assign Coef[802] = 'hE6214FE3ADDEF668E733FF1B7DED9C;
assign Coef[803] = 'hE2ABEFEF99D9C068E631FF3B7DE79C;
assign Coef[804] = 'hE72D6FE5ADDC0669EC31DF2B7D45DC;
assign Coef[805] = 'hE62F1FE7ABD88668E731DF3B7DD3DC;
assign Coef[806] = 'hD643621CF067355CEBBECBCBFD2C11;
assign Coef[807] = 'hDE117314B02615D2DBFCD9CFA90817;
assign Coef[808] = 'h1A535357A4241290DBFFDDC9920417;
assign Coef[809] = 'h12517217BC2010DADAFED9CBAB0A13;
assign Coef[810] = 'h76356B55FE20B9587ABECDCBABBB63;
assign Coef[811] = 'h5C306FB5A57293386932AB5DBBE9D2;
assign Coef[812] = 'h542A6DB6A53B9270E7A2AF1D3FE9F6;
assign Coef[813] = 'h64AA2DB0657C92686C2AAB1D7FE9E6;
assign Coef[814] = 'h64AA2FB5C57892686C2AA30D3FE1E6;
assign Coef[815] = 'hE66A4BB3451C83496C2EA71D2E41E6;
assign Coef[816] = 'hC76A4F93C53C8549FCAEAA9D6E4BCE;
assign Coef[817] = 'hC64A433BC1B91549FC8FAF9D644164;
assign Coef[818] = 'hD248456E8CB3F551F7D4A99B7CAD02;
assign Coef[819] = 'h50D2656EA8913D55F3D4ADDB799C10;
assign Coef[820] = 'hD070416E98F83DD1D0D58DCF599015;
assign Coef[821] = 'h5064707ED8F235DBD49ECDCB5D0A17;
assign Coef[822] = 'hC340772FB8B235DBD1D68DDBEB0C13;
assign Coef[823] = 'hD271D522E4E235D091F4CDC9F34853;
assign Coef[824] = 'hE2225483B570B1D0D0BCCF1BF9C05A;
assign Coef[825] = 'h42694FA39173B570F53ACFB979EBDE;
assign Coef[826] = 'hE2285DEF85DA9969F033CFBB7DE59E;
assign Coef[827] = 'hD308ECEFE1DB8768E463CFBB75FB1E;
assign Coef[828] = 'h4269AFADA5DAC669E423CF3B7DF5DE;
assign Coef[829] = 'hE22D6FEFADD8C769E621EF3B7DD5DC;
assign Coef[830] = 'hE62DE7EDADD8D768E4B17F29FDE5FE;
assign Coef[831] = 'h63275EEFC5D88628E4B1DF2BFD45DC;
assign Coef[832] = 'hF00369DD28063150623C8BCBA92571;
assign Coef[833] = 'hD011E354B2265154DBDA1B4BA20C12;
assign Coef[834] = 'h9A135217E42417D0D3FFDBCF820475;
assign Coef[835] = 'hE2537257B22630DAD8DED9CD8B0A43;
assign Coef[836] = 'hB6336EB5FA26BB5C78BECDCFABBF73;
assign Coef[837] = 'h54F26FB4C431937063328B1DBFE9C6;
assign Coef[838] = 'hDC126FB6853B9760E766AF9D7F6DC6;
assign Coef[839] = 'hD4220FB4C53B93286C22AF1D6FEDE6;
assign Coef[840] = 'h74AA0FA5455A8268642B230D6FE5E6;
assign Coef[841] = 'hEC6A0FB3C51A87497C2EA30F6E41E6;
assign Coef[842] = 'hC7424F83C5388349FC0DAA9F6E45CE;
assign Coef[843] = 'hDE4A43FBC59925496C85AF8F744184;
assign Coef[844] = 'hD842656EC09BB561F385AD9B79AC02;
assign Coef[845] = 'hD1D2656E1AB23DD5D3D4ADDB799401;
assign Coef[846] = 'hD042676E98B03DC3D0958DCB793017;
assign Coef[847] = 'hD640633FCABA394FD8972D8B0B4A17;
assign Coef[848] = 'hC350677ED2F235D3D1C68D8BE90E13;
assign Coef[849] = 'hDB5A752EE0F437D1D8F58DE9FB4857;
assign Coef[850] = 'hC6525D8AD9D0B1D0F0BFED2BFBE7DD;
assign Coef[851] = 'h404A6FA8F176B770F5BFCFBB79EBDE;
assign Coef[852] = 'hE2683CAA9DC27728E021CF2A79EFDE;
assign Coef[853] = 'hE2587BAF81DBE760E403EF2B7D699E;
assign Coef[854] = 'hE638BFAEC5DFE768E4214F2BFD6D9E;
assign Coef[855] = 'hE3ACAFEEEDDEE720E601EF3B7DF5DC;
assign Coef[856] = 'hE63DBFEDC9D8C768E401FF2B7D61DC;
assign Coef[857] = 'h473FFFADC5D9C728E401DF3FFDC5DE;
assign Coef[858] = 'hF2096A5D08C63D74F13B8B8BF36994;
assign Coef[859] = 'hB2516A55B0661756D3BA9B4B8A2E01;
assign Coef[860] = 'hB2537255B82513D2CAFFD94BD20C01;
assign Coef[861] = 'hB21372179A243FDED29CD9CD8B0343;
assign Coef[862] = 'h33016F15FC603F5CF8BE89CDAB8B02;
assign Coef[863] = 'h5C324F34C432937073328B19BBE0E2;
assign Coef[864] = 'hDC72DDB4457B9370EBE2AFBD7FECC6;
assign Coef[865] = 'h54328DB0455D9370EC20AB2975EDE6;
assign Coef[866] = 'hD4A80FA4457E8260E461AE0D7FE5E6;
assign Coef[867] = 'hFD220FB3451A87497C2EAE9F7E41E6;
assign Coef[868] = 'hE76A0F3BD5088549EC8FA98F2E05E6;
assign Coef[869] = 'hD6420BAAC5992741F48DAD9E7E4026;
assign Coef[870] = 'h5042416EB4933551D485A98B6D4802;
assign Coef[871] = 'hD0E0616EBCA33DF7F1D4ADCB799C01;
assign Coef[872] = 'h5460697EFAE03D46F095ADEBEB5175;
assign Coef[873] = 'hF622223BDAEA3D4FD09D2DCE1B4AB7;
assign Coef[874] = 'hC342437FDAE635CBD9C68D9B834E43;
assign Coef[875] = 'hD252F578DCC037D090DF8DBBE34457;
assign Coef[876] = 'hC270D782D1E027E0D09CEF3FFBE2D8;
assign Coef[877] = 'h42503F89D1C2BFE8E1A3CDBA79728D;
assign Coef[878] = 'hD4588DA8DDC28764C083EDAB7969CC;
assign Coef[879] = 'hF64CBBAEC9DAE760E501EFAB796CCC;
assign Coef[880] = 'hD238BDE885CE6764E501CF2B7D6D8C;
assign Coef[881] = 'hF62CAFEECDD8E764E401EF3B79F59C;
assign Coef[882] = 'hD63CAFECC1DB4728E4A1EF3B7D69CE;
assign Coef[883] = 'hD73EB5EB45D847A0E401FF2B7D55BC;
assign Coef[884] = 'hF008EBE808CEBF74E81D0A0ED905D0;
assign Coef[885] = 'hB211631590471B17D3FE8948C22C40;
assign Coef[886] = 'hBA13721FD26416D2D3BB59C9820643;
assign Coef[887] = 'hB6536A17FA2634D2F2BDD9C9922E21;
assign Coef[888] = 'hB3324F17DA6533DAF8BC899CA3ABA0;
assign Coef[889] = 'h1C528F96C40693D1F3A68BBDA3AD62;
assign Coef[890] = 'h5C525FB2842F97B1F3E0AB9DF2EC06;
assign Coef[891] = 'h5C30ADB4CC1F8320E461AF3DA764E6;
assign Coef[892] = 'hDC380DB4455E8231E4632B2D2EA5C6;
assign Coef[893] = 'hD4620FB3C5588349FC2CAB1F3F45C4;
assign Coef[894] = 'hD7020F9BD5188749FC2F2B862621A6;
assign Coef[895] = 'hD602033BC19A1743D48DAF8F744504;
assign Coef[896] = 'hD07A616E8E83BD73F584A98B790400;
assign Coef[897] = 'h00F0616E12823D67F094A99AC19C01;
assign Coef[898] = 'h7020E16EDAE2387750D48D8F499225;
assign Coef[899] = 'h7600633EDAF23C53D09D2D8B434E06;
assign Coef[900] = 'hB340626EDAE23DC3D18E888A830E01;
assign Coef[901] = 'h9652F30F58E03792D9F78D8AC34455;
assign Coef[902] = 'h5612F018D4C626F2D189EDADE54A2D;
assign Coef[903] = 'h6278B318D1EBA7E2D503CF282D6CCE;
assign Coef[904] = 'h5078AB6EC0C2A7E1F541CD2B516C85;
assign Coef[905] = 'h5628BFAC45C2E764E441CFAB7D6984;
assign Coef[906] = 'hF268BDAC05DF67A0E5036D297D698D;
assign Coef[907] = 'h7618BFECCDDFE76064006DABF9D5C5;
assign Coef[908] = 'hD638B5AECDD847A4E481EF2B7D65EC;
assign Coef[909] = 'hD63EBDEC4DD9C7A4E401CF2BF945ED;
assign Coef[910] = 'hB43A2E380E452F40A919880ED101A1;
assign Coef[911] = 'h3A50AE1398271F928BBBDA891B2C80;
assign Coef[912] = 'h93135201DA2537D0C2FBD9DE920623;
assign Coef[913] = 'hA2524A15DA273756FA9E48DCA20F22;
assign Coef[914] = 'h23326E17DE34B252F8BEC9DCAB0F20;
assign Coef[915] = 'h59125FB2841793B1FBFC8BBCBB8C50;
assign Coef[916] = 'h5C509FB2845793F1FBE78FBC2AEC02;
assign Coef[917] = 'h5D309FB0445382B1E422AA292A28E6;
assign Coef[918] = 'hDD1A8DB0445D82B1EE6F2E0C37A5E4;
assign Coef[919] = 'h5D6A8FF1C51A8741EC2FAB1E3605E6;
assign Coef[920] = 'hF5680F3BD51D0741F6AFAB967607A6;
assign Coef[921] = 'h56400379D61C0647EC8FAB9E2E0424;
assign Coef[922] = 'hD04A616CC2813D67F184A98A692E01;
assign Coef[923] = 'h10E0696EBA903D77DB142D8E819121;
assign Coef[924] = 'h7428615C5AC03877D2948D4E91B377;
assign Coef[925] = 'h3430A23C9A243E47D89CA98E8352E7;
assign Coef[926] = 'hB342603F9AA63CD7F88F888A032E03;
assign Coef[927] = 'hB210B178D0E316B7D49D898C964425;
assign Coef[928] = 'h1650D168D066B6D6D43DEBAAC52624;
assign Coef[929] = 'h3148093000E3B7B3F50DCDA8956C42;
assign Coef[930] = 'h3168A56C48C6EFE5E100EB2B41EC83;
assign Coef[931] = 'hF218AF6C82DAE7616700ED2B39FD06;
assign Coef[932] = 'h51789FA800EAE731E5406F2961EC24;
assign Coef[933] = 'h70389DEC80D8E76565006D2B796D65;
assign Coef[934] = 'h753CBDECCDDCC7A1E5006F297D6CE4;
assign Coef[935] = 'h963C9DAC40D967B4E601CF3B795C6D;
assign Coef[936] = 'h62E20CF84C95C805D39B810AF30CE1;
assign Coef[937] = 'h2A186A53AA673104B3F9C014562601;
assign Coef[938] = 'hBE7872219A241597C2BBD85A120601;
assign Coef[939] = 'hA7026E01DA643503FEBFD8CCD62260;
assign Coef[940] = 'hA0224E515874B616F83E8294828342;
assign Coef[941] = 'h09125E9A0C1437A1E2200A9CAB8560;
assign Coef[942] = 'h9952DDB2C49113B1DA640BBC326C66;
assign Coef[943] = 'hDD101DB0C47587B173E02A3C722C06;
assign Coef[944] = 'h5D109FB0041F83F1666BAB2C3FA0E6;
assign Coef[945] = 'h5D0A9F80851D82C17EAF2B963605A6;
assign Coef[946] = 'h4C4A0F31D55D27415EEFAF963625C6;
assign Coef[947] = 'h5440E33256D92467548DAC86044600;
assign Coef[948] = 'h1162E17A16832D277384A99A632701;
assign Coef[949] = 'h3080656E2A90BC7752148DFED99361;
assign Coef[950] = 'h3030E5587AE43E26D01C8DAE83B271;
assign Coef[951] = 'h35302E309A643E26518F4C029346A7;
assign Coef[952] = 'h2502425FDAA23CC3D18E088E470A23;
assign Coef[953] = 'h3010740892657E9190FDC80A064207;
assign Coef[954] = 'h1230B608B242B6A799094A3E45E642;
assign Coef[955] = 'h55788CB00263F72193618CAA35EC47;
assign Coef[956] = 'h711025E826C6BD2505010C282DEC67;
assign Coef[957] = 'h1270B56A2E5BE7656502CCA8696024;
assign Coef[958] = 'h1138B5A804EF7F25ED036F2A0C6504;
assign Coef[959] = 'hD178AD6CA8DAE72564006D2F69EDB7;
assign Coef[960] = 'h5728BDE004D946B44F40672A296845;
assign Coef[961] = 'h1C3C95AC6CC9E7B46401EF3B7D5475;
assign Coef[962] = 'hF0682CB886376325F81B038AEAAD71;
assign Coef[963] = 'h3842AA3B305601849C9B8198446C00;
assign Coef[964] = 'h163232119A2443829ABB5A544E0202;
assign Coef[965] = 'h2F142A63FB742600BC9BC0CE9E0672;
assign Coef[966] = 'hAE264A935A0497C0B2BA8C92C6A3A2;
assign Coef[967] = 'h9D525D020CA116E1C2EE89BE530C36;
assign Coef[968] = 'h9D121D920C31B791DB620B98AB2442;
assign Coef[969] = 'h981815A0845787B16BEE8B35380422;
assign Coef[970] = 'hDC521FA2441E86E1EE6EAEBD68E472;
assign Coef[971] = 'h7D129FB2455D03C1CC2A2F1F362064;
assign Coef[972] = 'h6D6207B0151E6447D62E2A167E0322;
assign Coef[973] = 'h750A832056902F674683AF167E0300;
assign Coef[974] = 'h0132617A2E936D67D2028BBAE99621;
assign Coef[975] = 'h20E2C92C7A8238675114097EC9B671;
assign Coef[976] = 'h2438801832027C26D01009E89196B3;
assign Coef[977] = 'h301A84A252302E2650AB858C83D2F3;
assign Coef[978] = 'hB142011B3A223D47908E888A0F8E23;
assign Coef[979] = 'h3918F00818E7368798AD091C462E33;
assign Coef[980] = 'hB05892821AE335A7800B812C2E4603;
assign Coef[981] = 'h98121D680E734707844605BA8DECC2;
assign Coef[982] = 'h157829486EC0FFA7CC068FBADDE863;
assign Coef[983] = 'h7C4E856804FB6FA54742092E09E866;
assign Coef[984] = 'h1D7895A820DB67A564068FB9497D21;
assign Coef[985] = 'h0138ADEEECFB6E2564000F2F79ED35;
assign Coef[986] = 'h503895AC48DD43B464400F2B6DCD77;
assign Coef[987] = 'h1C38BDA840D944B46600CF2B795137;
assign Coef[988] = 'hE00829E800DF69C1460E8718A10E11;
assign Coef[989] = 'hA14A22E13027CD068E9F80901C2EC2;
assign Coef[990] = 'h1B0BF6791A350B8687B9CB90560691;
assign Coef[991] = 'hAB034E03BA21CC470E3C809876A3A6;
assign Coef[992] = 'h2D2AAA13125681468E9F881AD6A7A3;
assign Coef[993] = 'h1932DD12543136C092EC809CE38887;
assign Coef[994] = 'h19125592245396819A6A0B987BAC32;
assign Coef[995] = 'h1912B5B684DFC2B1DBA80F38612422;
assign Coef[996] = 'hCC10B5A04404A7F5C76E8B3F7F0406;
assign Coef[997] = 'h0D2A17E2C45C0643DE2CAF3F570606;
assign Coef[998] = 'h5D2A8768DF1C25C3CCAEAB961E4744;
assign Coef[999] = 'h542201E82E4C45C346A48E362D2722;
assign Coef[1000] = 'hF06861DAB634FD67730009B6839371;
assign Coef[1001] = 'h20B2EC5C3E84B867701489FAD9D773;
assign Coef[1002] = 'h2430417032B62C06481C0D6C9392D1;
assign Coef[1003] = 'h24226C905A282E62802B060843F2E5;
assign Coef[1004] = 'h214060767A236D47910D19925A8E00;
assign Coef[1005] = 'h751074B2F82E56871EE30B2C1B4257;
assign Coef[1006] = 'hBE12B0D052776F861EABC0288FAE01;
assign Coef[1007] = 'h616011E11A67E7A21C278D28C44CC2;
assign Coef[1008] = 'hC568D86864D76D213C408D3C19DC75;
assign Coef[1009] = 'h416895CA0EEBEF6344448BBC09F835;
assign Coef[1010] = 'h111885CA6CFEC5775C008E29E9EC36;
assign Coef[1011] = 'hD4288D6800DD6D3444008F2CB9F837;
assign Coef[1012] = 'h5428ADE86CDBCEA44C000FAB29C905;
assign Coef[1013] = 'h1C38B5A864D863F445404FBF99CC77;
assign Coef[1014] = 'hA428256A2097C9078B1E810280CD11;
assign Coef[1015] = 'hE051304311978FA79E1D1098962A83;
assign Coef[1016] = 'h8A01EA72778C6A878EBD5010548792;
assign Coef[1017] = 'h2B00AEA7333C23468E2B1012462BAA;
assign Coef[1018] = 'h2F2AFED16BB503548C0E86103E83EB;
assign Coef[1019] = 'h8912F0020E0407F112AE89AED22662;
assign Coef[1020] = 'h8972D55A3CE517D198CE0E18D16400;
assign Coef[1021] = 'h9C52D5A464D527D19A648F19120C16;
assign Coef[1022] = 'h9812D1B2257D0791D0E28A1C5C0402;
assign Coef[1023] = 'hED1AD5664D0E06C14F6CAE3D0E07E6;
assign Coef[1024] = 'hCD52319A559E05C744ACAE8C360A02;
assign Coef[1025] = 'hF432AC7C638F4F6262AA8A1A5507C0;
assign Coef[1026] = 'h2060AD7C3A86AD475202891E9B8761;
assign Coef[1027] = 'hA0AAECAC7ED5FC679A12882A99F7F3;
assign Coef[1028] = 'hA40AC8807A26AF4668140D7CCBD293;
assign Coef[1029] = 'h240380B41B6C2A23080E401F97B790;
assign Coef[1030] = 'h210020441A46AD0218040492941EC1;
assign Coef[1031] = 'hA418F0D852F7A0831CAD4C3A4C2EE1;
assign Coef[1032] = 'h380AA07CDD26E1060EAF810A162A82;
assign Coef[1033] = 'h00323C7262F7C407866609A8ED2C83;
assign Coef[1034] = 'h854089346856EDA71E0005A849DDC7;
assign Coef[1035] = 'h081888F82076E5661D0605A8896976;
assign Coef[1036] = 'h4C3A9DAE207B85251D4401AF8DE857;
assign Coef[1037] = 'hC978CDA468DE44A569628F2BE9FDF7;
assign Coef[1038] = 'h1460FDB86CDB47F550208FBDE9FDB5;
assign Coef[1039] = 'h1C309DECE4C54BA04A600F3DD9DC35;
assign Coef[1040] = 'h80686C32245DED91167B048E5278D4;
assign Coef[1041] = 'hA80B3AC82B6E2F17941B108AA62218;
assign Coef[1042] = 'h0A61F24B7F8D43818E9F12C8460A8C;
assign Coef[1043] = 'h2529A6539BD5AD4A948B92922E278C;
assign Coef[1044] = 'h6F239283790622C69E2F949414A3CC;
assign Coef[1045] = 'h081250C21F2513908AAE0A99520662;
assign Coef[1046] = 'h0D53545A349625D2836E899AD25201;
assign Coef[1047] = 'h8859319AE45507919B6C8E80633E50;
assign Coef[1048] = 'h491BB1A2E4AF83A1C2E207BC176452;
assign Coef[1049] = 'h4C381560572C2180CEE6B4046C4240;
assign Coef[1050] = 'hCD421F244FED264756A8120C2C07C4;
assign Coef[1051] = 'h4C4350383B256E474E621C0C7C8325;
assign Coef[1052] = 'hA0AA897C3E0EAD064A0E81F2F9B631;
assign Coef[1053] = 'h21EBC85A2206AC260A1C815DB1F3F1;
assign Coef[1054] = 'hA0214CDC372CAA3648121CC09BD3D7;
assign Coef[1055] = 'hA021E8F65B65AE2600055418DFEEFD;
assign Coef[1056] = 'hE003181D1222AC42080D141A87DAC2;
assign Coef[1057] = 'h040A2054F2A64C0616EB1A1AD66E83;
assign Coef[1058] = 'h443BBC632FE60CA39C0F13AAAC7EA0;
assign Coef[1059] = 'h24031C307AE32D0300431320EC2E10;
assign Coef[1060] = 'h68787C8646FCCA2750261998CCCD74;
assign Coef[1061] = 'h2548B1E820F3EF3354000DB349C855;
assign Coef[1062] = 'hDC71BD9E6CD06DF14840073799EDF7;
assign Coef[1063] = 'h4D39BCBC6CF764A5CA400FBBF9DC17;
assign Coef[1064] = 'h086BEDA2A461C1B1422203AD89E8F5;
assign Coef[1065] = 'h5C317D8C40CAC6B448440563F9D0B5;
assign Coef[1066] = 'hB441247A04D72B0292278592260457;
assign Coef[1067] = 'h84C9F82B37BDA94A92C6971844B699;
assign Coef[1068] = 'h25093019BBE40B171E0B1458DCB689;
assign Coef[1069] = 'h416BAC79191C0056A62B10168657CC;
assign Coef[1070] = 'h2C6ADCF3F36441278E2F94989E12BE;
assign Coef[1071] = 'h895374D333D593919A2C960C3A064C;
assign Coef[1072] = 'h895B545A943107919A42965A6A2407;
assign Coef[1073] = 'h590210BAEC43C7909BEF8BFF3A0050;
assign Coef[1074] = 'h581BD522E49FC4919AE20FBE162402;
assign Coef[1075] = 'h791835656F1FC6D34C4B9F3F2E2004;
assign Coef[1076] = 'hDD4A94F8671C47474E8F3E0B6E0600;
assign Coef[1077] = 'hE92A48E33FBC8C02462295120EA715;
assign Coef[1078] = 'hE1E8E5C64A0DAF23B2268038EBBFD1;
assign Coef[1079] = 'h21EA484FB38EA92E881C10F2C993B1;
assign Coef[1080] = 'h25B8688E7FAAE826200209F8C2F79D;
assign Coef[1081] = 'h64498819130E804A9C2F940C8CBFCA;
assign Coef[1082] = 'hA17800A213EE8C1E25291042AA4EE6;
assign Coef[1083] = 'hED1924533B7A47031CEF92300E469C;
assign Coef[1084] = 'h447A0C30673F0B020461D3AC566C64;
assign Coef[1085] = 'h6D09381AE384CC161FAB812BFEFCF6;
assign Coef[1086] = 'hAC3964D40AD157E1122689A8D9D815;
assign Coef[1087] = 'h8D6A1844E0C766B340408FBFB96973;
assign Coef[1088] = 'h591B44C459DF60B518E68FECBBED37;
assign Coef[1089] = 'h89789474A0E0B995D1420BEB895D93;
assign Coef[1090] = 'h0819DC442C6A72B349460729D99473;
assign Coef[1091] = 'h183190DA80F9F0B4D0628F3FF9DC73;
assign Coef[1092] = 'h882D307B5BDD895EB9221402125621;
assign Coef[1093] = 'hA14B003915CD0BDA1026128274170A;
assign Coef[1094] = 'hA50BB26B0F942E5B9E09109866D48C;
assign Coef[1095] = 'hE40D6623DBDC85DB260B10946C678C;
assign Coef[1096] = 'h0C4B10F1530C00D28409D29F5697EE;
assign Coef[1097] = 'h2913544F106C6B12838E14FA96768E;
assign Coef[1098] = 'h8553501A62276C921AE490C27C0441;
assign Coef[1099] = 'h1A05B83E34B7079393C60E3876344A;
assign Coef[1100] = 'hCD1390467CDB60D982EF06DC6C6646;
assign Coef[1101] = 'hCD1B11E80DDC43DC44EB361C462C43;
assign Coef[1102] = 'h5C3E54694F9C0BDF0ECFBA16740208;
assign Coef[1103] = 'h64336851139CC162564F94763965A5;
assign Coef[1104] = 'h60F86C7F720C6B5EEA00842C29F773;
assign Coef[1105] = 'h24B34C042B04A83E2B100062C1FFF3;
assign Coef[1106] = 'hA5698CB47F3DA22A2E180020A2BFED;
assign Coef[1107] = 'h6419A8A95F2ACD36BC08821096F6CE;
assign Coef[1108] = 'hC00DAC1B1B2E8A3A2D6D91F2BEEBC9;
assign Coef[1109] = 'h640D3C8E93AAC8BB1C6F90406E0C8A;
assign Coef[1110] = 'h7C7BDCAB27D7501A14A29092246EAE;
assign Coef[1111] = 'h611BB023BB6143B2264612ACAC6822;
assign Coef[1112] = 'hA469080C74F6E216080E84EC528CC5;
assign Coef[1113] = 'h4937848044F3FDBA80268CA8ABADBD;
assign Coef[1114] = 'h08315D3428E253B48A660EE99B8817;
assign Coef[1115] = 'h8839D4C24475D89010220DFBA9CD37;
assign Coef[1116] = 'h4839146464F353315360856E69AC57;
assign Coef[1117] = 'h0C799CECE4F6EBB0C2628F6AB9DC77;
assign Coef[1118] = 'hB0AA643B420DE91A38461080E264DE;
assign Coef[1119] = 'hAF69C7A33F7D485ABD18B412B88709;
assign Coef[1120] = 'h863F142F3B2E891E0F62B29B761F08;
assign Coef[1121] = 'hEA2B16F9575E829AA70DA2444EB4BE;
assign Coef[1122] = 'hEF734AA31772635A3C6BD4164E5629;
assign Coef[1123] = 'h8A41205364F462928AC815D2562805;
assign Coef[1124] = 'h8B1D301A5F97E3920A4006A070940F;
assign Coef[1125] = 'hCF7B15622CB5679093EB90EE541C54;
assign Coef[1126] = 'h5A3850214C9D479095EA19124C0A60;
assign Coef[1127] = 'h7F1895BBDF9403D144E93B302E24E6;
assign Coef[1128] = 'h586B1FA3F35E46DA962B14A254650D;
assign Coef[1129] = 'hE888FFA907560A886C0312222E07C2;
assign Coef[1130] = 'hE4A96C6C6A56D96E295823BED9B776;
assign Coef[1131] = 'hA0EB08C63A0EA03E221293ECAB9989;
assign Coef[1132] = 'hA48B88C4626699ACA60AA2A6919FC8;
assign Coef[1133] = 'hA0083895371D6C4A356986E43F7DEF;
assign Coef[1134] = 'h655B099B3234AB8E3D4C4406355E8E;
assign Coef[1135] = 'h650AA679336D891B1441D364B685C4;
assign Coef[1136] = 'hE01138343A12F7183E2890AB460FC0;
assign Coef[1137] = 'h204818574DBFE12A2664BD1DA85E26;
assign Coef[1138] = 'h806BA8242867697C994613E0BBDC54;
assign Coef[1139] = 'h80138CB612016F74D8468DB9CAF673;
assign Coef[1140] = 'h8539E89C48BFFB3029060FEADBEE77;
assign Coef[1141] = 'h8DF9C08CACBE51FCC1240F6EB9DCF3;
assign Coef[1142] = 'h1419C0307843589C9A00877AA9D457;
assign Coef[1143] = 'h1939DC8CCC675194DA4283E8ABECB3;
assign Coef[1144] = 'h8B8A23F13A2CE9E9020C2022407EC5;
assign Coef[1145] = 'hAA0B22AB02BCC24E2447D112041448;
assign Coef[1146] = 'h8B3B261952D4C386AE13329234A74B;
assign Coef[1147] = 'h6B0B16ED19DDC0228E091696242FB8;
assign Coef[1148] = 'hBE6B13D9732D6ACABE29D000348DEF;
assign Coef[1149] = 'h9B5A965B794DC2821AA7949ED4048D;
assign Coef[1150] = 'h991B7003F1A772D397EAD44CD8340D;
assign Coef[1151] = 'h9A49162A2D0577F409EB107A020213;
assign Coef[1152] = 'hBF4BB24B308583822AAF54B234180A;
assign Coef[1153] = 'h8D0912B347BF61C0CEEFB6B4460A2C;
assign Coef[1154] = 'h5F109ACA5E0F44E21F6DB6846C448C;
assign Coef[1155] = 'hD73828395693436D2E43B0061CBE9D;
assign Coef[1156] = 'hE4C9AC4D620C5B2EB116000C39D568;
assign Coef[1157] = 'h60A988C63A40C86A290022C5C3BF8D;
assign Coef[1158] = 'hE3A92C811C56E0AE081EE6ACFD7FF8;
assign Coef[1159] = 'hEFAB2090B3ACC10E3C27262016F6EC;
assign Coef[1160] = 'hE6EA8AD2129EE128360020D70466ED;
assign Coef[1161] = 'h72392CB927EE4B16BC6FA6A4BE24E4;
assign Coef[1162] = 'hE3393216D21BB13A8D0735A69E448C;
assign Coef[1163] = 'hCD8B22B45A6C2986B828B164CBEE42;
assign Coef[1164] = 'hA55B18224443F1725924471D19D499;
assign Coef[1165] = 'h91A3D86074D773303024CC4D6BDC57;
assign Coef[1166] = 'h107961D632C0F9D08A6605689BFED1;
assign Coef[1167] = 'h9DB954E63C70D8B008780768BBEEF7;
assign Coef[1168] = 'h895BC4FC4CEDF81409568F7D9970F5;
assign Coef[1169] = 'h0D185C484CE4DBB0183603E9B9F0F7;
assign Coef[1170] = 'hBDCC423D7CFFEC5AAD030590443E1F;
assign Coef[1171] = 'hAA0DA71F312F255F360B11825C9729;
assign Coef[1172] = 'hC0A9037B1A948A673E179033645284;
assign Coef[1173] = 'hF6AE83D71F5FC044B62BB3176E219C;
assign Coef[1174] = 'h87AAA62BD3D440D2FEA07240262E88;
assign Coef[1175] = 'hFF4B306BDFA54892A40D3047D4140C;
assign Coef[1176] = 'hCE5F5213150751C39D7550B04E0219;
assign Coef[1177] = 'hF31EB23627A550F492EFD7925A0408;
assign Coef[1178] = 'hDE0C32FBA5965990886B9260060244;
assign Coef[1179] = 'h5C0892A2C5AD5A9946C19033040E1C;
assign Coef[1180] = 'hF31A3F698F2E41D0D76F106522011C;
assign Coef[1181] = 'h79688355CB1D6A7CEF011477604C58;
assign Coef[1182] = 'hA1A8A98F463CD93E623AB5F16BB5DD;
assign Coef[1183] = 'hE1AC0D0D43FDE86E301084A5D3F5F6;
assign Coef[1184] = 'hA4A9EFC45B04EA4CEB1E66639DCFA8;
assign Coef[1185] = 'h7529AAA1075EA9687E2800E7B6A5E8;
assign Coef[1186] = 'h71A90F951BB74E3E2E0CA290F093C8;
assign Coef[1187] = 'hFDCE3AEA152668BAADD9F3D0CE409A;
assign Coef[1188] = 'hFE0B2B554059D008BFE202A72237D9;
assign Coef[1189] = 'hE909021B736CC352910891C13FDE71;
assign Coef[1190] = 'hC9BD09960A75DA94985685AFD9E856;
assign Coef[1191] = 'h9D31FD4576E4D8D6A17606F6D3DD33;
assign Coef[1192] = 'h84B9ED843075F0F011FE83E989F651;
assign Coef[1193] = 'h8899654430F7F8B10956836BB35873;
assign Coef[1194] = 'h0199DD7E4C677394C9F2877FBBF957;
assign Coef[1195] = 'h083BD1DC64A47AB4D1361FECE96C17;
assign Coef[1196] = 'h124AB563E4D7D8CC229EB012207660;
assign Coef[1197] = 'hF04E237B5A97EDCC3E5334A4243F89;
assign Coef[1198] = 'hF2EF773BDFDC49C6060FA4D2658213;
assign Coef[1199] = 'h6FFF033A3F0DEE62342B320426E78D;
assign Coef[1200] = 'h7A4DA7E90F8D29CA86AFF032442CA8;
assign Coef[1201] = 'h9A2EB049245E409AAEA942D0362A05;
assign Coef[1202] = 'hDF5BF45B31862782BEC3D2475E0E2B;
assign Coef[1203] = 'hDB4F16C3158F47D01BEB85736C2E0A;
assign Coef[1204] = 'hDE199178BF2544C496E3F7C41C2C4A;
assign Coef[1205] = 'hDE3B77070D8C48F184C316C07E2C1B;
assign Coef[1206] = 'hDC0A128ADDCCC220D09334343E06CE;
assign Coef[1207] = 'hDEB9872D691ECA4ABE4F95245ACC0B;
assign Coef[1208] = 'hF4AD2D85023FCA2FEE4FA1A6AA9537;
assign Coef[1209] = 'hE5EBEFA963B4FB2E32162530DBF0C4;
assign Coef[1210] = 'h71AB8D3BD11EF92C201BD210A9F3E4;
assign Coef[1211] = 'hF5EB6703736E4A0E053B304C0FD34F;
assign Coef[1212] = 'hE72B09F763940A0E361BB080AE97AC;
assign Coef[1213] = 'hEAE9A93432A5613A58EAC3D3F264B5;
assign Coef[1214] = 'hFE531B68016DC60E081B1719DC5C3C;
assign Coef[1215] = 'hA737D08E9E25E92410331368ADCC44;
assign Coef[1216] = 'hC30BD8546246C073D8FE8BD88394B6;
assign Coef[1217] = 'h492B59166AE63A0FDA7283F889CEF7;
assign Coef[1218] = 'h07FBC564A856F930905205EE89EE91;
assign Coef[1219] = 'h105944964874F1B2887AC76EEBEC73;
assign Coef[1220] = 'h901B74D424AD53B491748F6A99EA57;
assign Coef[1221] = 'h813BDCF424877E94E976476C81E4D1;
assign Coef[1222] = 'hC6C9F67202CEFB6AEF9225231FE400;
assign Coef[1223] = 'hA2BA036D3F1FCD1A7C4B7422646840;
assign Coef[1224] = 'hEEEE23791F37697F3F4FB4925C06AF;
assign Coef[1225] = 'hEB0A2639559ECA4EEC0772907E5068;
assign Coef[1226] = 'hFE0CB63BD78D60F0F60B330656338E;
assign Coef[1227] = 'hBF0A32092B844FB4328F95325E1ECC;
assign Coef[1228] = 'h125F90C375A54CD29DE3D2B50E0A1F;
assign Coef[1229] = 'hDF0AB262820F748885E330D93C4C0D;
assign Coef[1230] = 'h5A1B927A27D756C297CA5D55260E9D;
assign Coef[1231] = 'hEB1DB28B0D3C43705EEB16261C0D99;
assign Coef[1232] = 'hDB8FB5291CDE4728CFDB32B6040CCE;
assign Coef[1233] = 'hEC48A7A5C5DDCDF52D0665B4071D3E;
assign Coef[1234] = 'hE1288D6C764FD07E600A20E2DDB7B8;
assign Coef[1235] = 'h84A90DC40936E82C881EE2AB9BDF9C;
assign Coef[1236] = 'hC6AC2AD4511EC22C7A12E19C5F94EC;
assign Coef[1237] = 'hB4CAAFF49C6C495ECC6EA63B5A91BE;
assign Coef[1238] = 'hC42D4A7F5F0C8F03E417B68529FAFA;
assign Coef[1239] = 'h36D829B55C5ECA7A206EA2426FF04E;
assign Coef[1240] = 'hA2FBBB2B19844606901FE331F97A45;
assign Coef[1241] = 'h44C9EC9D1B65F3FABA5EF0EAD32ECF;
assign Coef[1242] = 'hB6394D8C88F5721EBB761DF981E8F2;
assign Coef[1243] = 'hBFF968946A75D0F48B1A0A6FAB4E11;
assign Coef[1244] = 'h01B95D4438F5F3D99972C5FE81B071;
assign Coef[1245] = 'h01F9DD4EE2E478941AF20D4FB9F675;
assign Coef[1246] = 'h981BD18628D6F3901B7E8769B9C873;
assign Coef[1247] = 'h88B9D0AC5CD5F0B0C9724FE9CBF811;
assign Coef[1248] = 'hB8EB473B821FFFCB4FE730643C7106;
assign Coef[1249] = 'hF4C93623573CFD96AF43520B6CB684;
assign Coef[1250] = 'hE3ACA77B549F635FF6EF70BE0606C2;
assign Coef[1251] = 'hC7EE01B547FD610E5E4B7597D40D8C;
assign Coef[1252] = 'h4AAA22A1B1C5446A1CC3F6824E428A;
assign Coef[1253] = 'h162F93DF1B8646E89DABD213542A8C;
assign Coef[1254] = 'hB81B23D92BE4C194ADEFD2D564410B;
assign Coef[1255] = 'h9A1B526816CF4D9A87C736C1000005;
assign Coef[1256] = 'hFF1F93687CA747DB97E7636D6C0C06;
assign Coef[1257] = 'h5F0883E1CF5E47DAC5AFF6756642CA;
assign Coef[1258] = 'h568A8FF2C41FE358E0EF382E65608A;
assign Coef[1259] = 'hECBA139306AFE96AE80BA79535262C;
assign Coef[1260] = 'hB1E8ACC97B76FB2C3A4EE0BE79DBDB;
assign Coef[1261] = 'hEDAFE9C7465FD90EE25EA008D5F5EE;
assign Coef[1262] = 'hB19B29254F2C6A3C2D1AA5F333C7DC;
assign Coef[1263] = 'h77AFAEFF2B5D46A8AD23616D19DFBA;
assign Coef[1264] = 'h112EADE74B1EF2BF7A8BC22ACF6BE4;
assign Coef[1265] = 'hA2582F08F16EEE2AE9FE322BED6B06;
assign Coef[1266] = 'hAE996E474147F77ECB8A65FF33BC3B;
assign Coef[1267] = 'hCE3B0997726C5056D2A655CAFBDEEB;
assign Coef[1268] = 'h02B9C1D60AE5FB13839E84EFA9ACF1;
assign Coef[1269] = 'hA1FBD14C8CA6799EAA7EC568939AF5;
assign Coef[1270] = 'hA0B9DDDC44A479B249F6C5C893A871;
assign Coef[1271] = 'h001BC9CE2E6579B4D8B2CFEB83E833;
assign Coef[1272] = 'h1DDBD45C3865FB9CAB52C77A9BB851;
assign Coef[1273] = 'h081BD446ACA67390D07EC77DD3F473;



assign   coef= Coef[addr];
endmodule