/*
date:2018/5/8
���ںţ�С��FPGA
���ں��ϡ���2Ƶ��FFTʵ��-verilogƪ2�������̽���
*/

module fw_sram_2 #(
  parameter WIDTH_A = 12
)
(
   input [WIDTH_A-1:0] addr,
   
   output[79:0]  coef

);

       

wire [79:0] Coef [0:119];
assign Coef[0] = 'h40C92A00B164044E689A;
assign Coef[1] = 'h00107F11504205020076;
assign Coef[2] = 'h2113C90CACEA232E28B7;
assign Coef[3] = 'h5D52B4E0509455C501C8;
assign Coef[4] = 'hDD206B6353135C990488;
assign Coef[5] = 'h3113FB526882061120FE;
assign Coef[6] = 'hC5F81BA193558D4DF146;
assign Coef[7] = 'hB1CD52B7B54CBD776F83;
assign Coef[8] = 'h6429F36BEA75C9AE295B;
assign Coef[9] = 'hE6EB00B7F57DDBEFCE00;
assign Coef[10] = 'h2306C94C2CC301220A5E;
assign Coef[11] = 'h1B30E440429054492608;
assign Coef[12] = 'h157FBCD4E54F529F8BFC;
assign Coef[13] = 'h66FB28D9ABD189E8A14E;
assign Coef[14] = 'h421052A4346120C26DC5;
assign Coef[15] = 'hD5A8EF09FB906DD9E915;
assign Coef[16] = 'h0DF4AE461BA24A9D8158;
assign Coef[17] = 'h14686E0CE4841D877D92;
assign Coef[18] = 'hF7CBADCF95469CC94A96;
assign Coef[19] = 'hDFB2227B1B9DFC787508;
assign Coef[20] = 'h092D6A0446B245821A62;
assign Coef[21] = 'h795F3E46A6261F6B0799;
assign Coef[22] = 'hC5B9E3B7BB46ADFF89E4;
assign Coef[23] = 'h18D736B6B54241D7CEF2;
assign Coef[24] = 'h3515AE4D1593E42081B9;
assign Coef[25] = 'h086ED9FCA46DBDFE79DE;
assign Coef[26] = 'hBFDFBDDCFCCF9E6F4AB0;
assign Coef[27] = 'h7B5AA9ADFD96DC0FD421;
assign Coef[28] = 'hEEEC56FA810D1B7C775F;
assign Coef[29] = 'h15C8CE45A144494EE95E;
assign Coef[30] = 'h68C9D4AA904429777C0B;
assign Coef[31] = 'hA1F80BA5FB4ACD4E89C7;
assign Coef[32] = 'h50883B0522E444436184;
assign Coef[33] = 'h33108A1438A201032BDC;
assign Coef[34] = 'hD6FE8FF4AF5DFAEAD184;
assign Coef[35] = 'hE6A95B07E3FFEC3EE9A6;
assign Coef[36] = 'h2949C914F46EB5DE7EBB;
assign Coef[37] = 'h9912BE725807355927DF;
assign Coef[38] = 'h65ECC91FECE3C7AE6B67;
assign Coef[39] = 'h6532EA195BB2C4230176;
assign Coef[40] = 'hDE6476FB47081BD0675D;
assign Coef[41] = 'h7D96FFED4D825649821E;
assign Coef[42] = 'h6FF88125E5C47D9D7481;
assign Coef[43] = 'hF95FBD56FD6F1FCB48BE;
assign Coef[44] = 'h251AFF4BD882444A807E;
assign Coef[45] = 'h35F3EA13335485C549E6;
assign Coef[46] = 'h7BFDB43BD4975DEFC4A1;
assign Coef[47] = 'hFFFE37D3D37F5BE9C69C;
assign Coef[48] = 'h64FF2657E7F369E6C6B1;
assign Coef[49] = 'h6FFEA76FF7C459DD4D4A;
assign Coef[50] = 'h62EF0A0CC7C63D5EEE12;
assign Coef[51] = 'h18406645E056578DEE88;
assign Coef[52] = 'hAECFCB4D8D4BAF7E7AFF;
assign Coef[53] = 'h54FA32A7B3440BCDFDC0;
assign Coef[54] = 'h77B46E435392E441F385;
assign Coef[55] = 'h00FD44ACF54415FE4663;
assign Coef[56] = 'hFB32EF784A9D9A19F408;
assign Coef[57] = 'h00581048F076090EEC26;
assign Coef[58] = 'h3707EE4B55931460867F;
assign Coef[59] = 'h5DE06E4102941601808C;
assign Coef[60] = 'h45606A0161D2458C0D44;
assign Coef[61] = 'hE3EF8F4DBFFFDD6C0956;
assign Coef[62] = 'h04CBCB1DE5D7878EE9A7;
assign Coef[63] = 'hB47F07B6B06F23357DF6;
assign Coef[64] = 'h6CA95AAF111D1EE36A73;
assign Coef[65] = 'h1520C6697A1041824DB0;
assign Coef[66] = 'h457D2A04F7722BE689D6;
assign Coef[67] = 'h62A9C81EC9A68FFE6CA3;
assign Coef[68] = 'h0506DE00E4E2440FFD8C;
assign Coef[69] = 'h23327BB35233CB2181F4;
assign Coef[70] = 'h9AB632F2523DAB85CFDD;
assign Coef[71] = 'h58F922B5D864B9FDC6C9;
assign Coef[72] = 'hCFFAF3F0F1CCDE5D7C82;
assign Coef[73] = 'h5BF077624235DFE98701;
assign Coef[74] = 'h191392415B30E411B1BE;
assign Coef[75] = 'h5DA1EF49EBD05D0DA9CF;
assign Coef[76] = 'h23339B0376F7E12349A7;
assign Coef[77] = 'hA5FB12BDFC47EDBE7E83;
assign Coef[78] = 'h01C907A7DAE66947C8C0;
assign Coef[79] = 'hEF9174FB1B38EFE183FE;
assign Coef[80] = 'hE8CF8006B46715D64EB0;
assign Coef[81] = 'h47A8C20543988D6D8146;
assign Coef[82] = 'hE0995BF3CC4F40E649FE;
assign Coef[83] = 'hC328EBA8EB84CDCE6146;
assign Coef[84] = 'h01A076C062C65D4EFCE0;
assign Coef[85] = 'h199EECCC2C82134B0290;
assign Coef[86] = 'h1B15F6E256924401877C;
assign Coef[87] = 'h1D880A45E2C245512CBE;
assign Coef[88] = 'hCEE94086E35DFBFEEEA0;
assign Coef[89] = 'h4DE8E56D6F99BFC9E441;
assign Coef[90] = 'h0400661147A074080648;
assign Coef[91] = 'h481854B452401082C4B8;
assign Coef[92] = 'h09EC2808E7D40956D9D4;
assign Coef[93] = 'h1306F1863029B4A21BFE;
assign Coef[94] = 'h02004A0CA0420012085E;
assign Coef[95] = 'h1548EE414044454001D4;
assign Coef[96] = 'hC9CC6245C5807DD07F5B;
assign Coef[97] = 'h48850EF317017931877E;
assign Coef[98] = 'h3CD73646F44623EF42B4;
assign Coef[99] = 'h9A0516F05631F261A57C;
assign Coef[100] = 'h052462446004454041F0;
assign Coef[101] = 'h1333FBB21233C42309E4;
assign Coef[102] = 'hA15A8137FAD6C2AB3CA7;
assign Coef[103] = 'h04C4244DE6C05588A22A;
assign Coef[104] = 'h29CDCC44E7C2610C8B5F;
assign Coef[105] = 'hBD1CECC94DC352090630;
assign Coef[106] = 'hFDFFA515E7F35FCAC6A1;
assign Coef[107] = 'h64EECF4DC99117EC0F4F;
assign Coef[108] = 'h4CF830ADED66DBFFF481;
assign Coef[109] = 'h4AB531311335EBC5CF47;
assign Coef[110] = 'hC4FADB1EEFFFEF7E78A6;
assign Coef[111] = 'h25608B0CDEC305E68944;
assign Coef[112] = 'h2117CB114DA2E626097F;
assign Coef[113] = 'h9907A82CAC42A74D67DB;
assign Coef[114] = 'h2116DA4468C25322299E;
assign Coef[115] = 'h5D10EE494AC055C8110C;
assign Coef[116] = 'hE5736F2B4FA98979811F;
assign Coef[117] = 'h1B1426275892420308DC;
assign Coef[118] = 'h18552284F43293A3C681;
assign Coef[119] = 'hDADC9DD4C8CCBBDD7C4F;



assign   coef= Coef[addr];
endmodule